VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO mp3_data_array_2
   CLASS BLOCK ;
   SIZE 893.635 BY 127.445 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  161.69 1.0375 161.825 1.1725 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  164.55 1.0375 164.685 1.1725 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  167.41 1.0375 167.545 1.1725 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  170.27 1.0375 170.405 1.1725 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  173.13 1.0375 173.265 1.1725 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  175.99 1.0375 176.125 1.1725 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.85 1.0375 178.985 1.1725 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  181.71 1.0375 181.845 1.1725 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  184.57 1.0375 184.705 1.1725 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  187.43 1.0375 187.565 1.1725 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  190.29 1.0375 190.425 1.1725 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  193.15 1.0375 193.285 1.1725 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  196.01 1.0375 196.145 1.1725 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  198.87 1.0375 199.005 1.1725 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  201.73 1.0375 201.865 1.1725 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  204.59 1.0375 204.725 1.1725 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  207.45 1.0375 207.585 1.1725 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  210.31 1.0375 210.445 1.1725 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  213.17 1.0375 213.305 1.1725 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  216.03 1.0375 216.165 1.1725 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  218.89 1.0375 219.025 1.1725 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  221.75 1.0375 221.885 1.1725 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  224.61 1.0375 224.745 1.1725 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  227.47 1.0375 227.605 1.1725 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  230.33 1.0375 230.465 1.1725 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  233.19 1.0375 233.325 1.1725 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  236.05 1.0375 236.185 1.1725 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  238.91 1.0375 239.045 1.1725 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  241.77 1.0375 241.905 1.1725 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  244.63 1.0375 244.765 1.1725 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  247.49 1.0375 247.625 1.1725 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  250.35 1.0375 250.485 1.1725 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  253.21 1.0375 253.345 1.1725 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  256.07 1.0375 256.205 1.1725 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  258.93 1.0375 259.065 1.1725 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  261.79 1.0375 261.925 1.1725 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  264.65 1.0375 264.785 1.1725 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  267.51 1.0375 267.645 1.1725 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  270.37 1.0375 270.505 1.1725 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  273.23 1.0375 273.365 1.1725 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  276.09 1.0375 276.225 1.1725 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  278.95 1.0375 279.085 1.1725 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  281.81 1.0375 281.945 1.1725 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  284.67 1.0375 284.805 1.1725 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  287.53 1.0375 287.665 1.1725 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  290.39 1.0375 290.525 1.1725 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  293.25 1.0375 293.385 1.1725 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  296.11 1.0375 296.245 1.1725 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  298.97 1.0375 299.105 1.1725 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  301.83 1.0375 301.965 1.1725 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  304.69 1.0375 304.825 1.1725 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  307.55 1.0375 307.685 1.1725 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  310.41 1.0375 310.545 1.1725 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  313.27 1.0375 313.405 1.1725 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  316.13 1.0375 316.265 1.1725 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  318.99 1.0375 319.125 1.1725 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  321.85 1.0375 321.985 1.1725 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  324.71 1.0375 324.845 1.1725 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  327.57 1.0375 327.705 1.1725 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  330.43 1.0375 330.565 1.1725 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  333.29 1.0375 333.425 1.1725 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  336.15 1.0375 336.285 1.1725 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  339.01 1.0375 339.145 1.1725 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  341.87 1.0375 342.005 1.1725 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  344.73 1.0375 344.865 1.1725 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  347.59 1.0375 347.725 1.1725 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  350.45 1.0375 350.585 1.1725 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  353.31 1.0375 353.445 1.1725 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  356.17 1.0375 356.305 1.1725 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  359.03 1.0375 359.165 1.1725 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  361.89 1.0375 362.025 1.1725 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  364.75 1.0375 364.885 1.1725 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  367.61 1.0375 367.745 1.1725 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  370.47 1.0375 370.605 1.1725 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  373.33 1.0375 373.465 1.1725 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  376.19 1.0375 376.325 1.1725 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  379.05 1.0375 379.185 1.1725 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  381.91 1.0375 382.045 1.1725 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  384.77 1.0375 384.905 1.1725 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  387.63 1.0375 387.765 1.1725 ;
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  390.49 1.0375 390.625 1.1725 ;
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  393.35 1.0375 393.485 1.1725 ;
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  396.21 1.0375 396.345 1.1725 ;
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  399.07 1.0375 399.205 1.1725 ;
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  401.93 1.0375 402.065 1.1725 ;
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  404.79 1.0375 404.925 1.1725 ;
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  407.65 1.0375 407.785 1.1725 ;
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  410.51 1.0375 410.645 1.1725 ;
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  413.37 1.0375 413.505 1.1725 ;
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  416.23 1.0375 416.365 1.1725 ;
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  419.09 1.0375 419.225 1.1725 ;
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  421.95 1.0375 422.085 1.1725 ;
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  424.81 1.0375 424.945 1.1725 ;
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  427.67 1.0375 427.805 1.1725 ;
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  430.53 1.0375 430.665 1.1725 ;
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  433.39 1.0375 433.525 1.1725 ;
      END
   END din0[95]
   PIN din0[96]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  436.25 1.0375 436.385 1.1725 ;
      END
   END din0[96]
   PIN din0[97]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  439.11 1.0375 439.245 1.1725 ;
      END
   END din0[97]
   PIN din0[98]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  441.97 1.0375 442.105 1.1725 ;
      END
   END din0[98]
   PIN din0[99]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  444.83 1.0375 444.965 1.1725 ;
      END
   END din0[99]
   PIN din0[100]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  447.69 1.0375 447.825 1.1725 ;
      END
   END din0[100]
   PIN din0[101]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  450.55 1.0375 450.685 1.1725 ;
      END
   END din0[101]
   PIN din0[102]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  453.41 1.0375 453.545 1.1725 ;
      END
   END din0[102]
   PIN din0[103]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  456.27 1.0375 456.405 1.1725 ;
      END
   END din0[103]
   PIN din0[104]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  459.13 1.0375 459.265 1.1725 ;
      END
   END din0[104]
   PIN din0[105]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  461.99 1.0375 462.125 1.1725 ;
      END
   END din0[105]
   PIN din0[106]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  464.85 1.0375 464.985 1.1725 ;
      END
   END din0[106]
   PIN din0[107]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  467.71 1.0375 467.845 1.1725 ;
      END
   END din0[107]
   PIN din0[108]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  470.57 1.0375 470.705 1.1725 ;
      END
   END din0[108]
   PIN din0[109]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  473.43 1.0375 473.565 1.1725 ;
      END
   END din0[109]
   PIN din0[110]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  476.29 1.0375 476.425 1.1725 ;
      END
   END din0[110]
   PIN din0[111]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  479.15 1.0375 479.285 1.1725 ;
      END
   END din0[111]
   PIN din0[112]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  482.01 1.0375 482.145 1.1725 ;
      END
   END din0[112]
   PIN din0[113]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  484.87 1.0375 485.005 1.1725 ;
      END
   END din0[113]
   PIN din0[114]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  487.73 1.0375 487.865 1.1725 ;
      END
   END din0[114]
   PIN din0[115]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  490.59 1.0375 490.725 1.1725 ;
      END
   END din0[115]
   PIN din0[116]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  493.45 1.0375 493.585 1.1725 ;
      END
   END din0[116]
   PIN din0[117]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  496.31 1.0375 496.445 1.1725 ;
      END
   END din0[117]
   PIN din0[118]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  499.17 1.0375 499.305 1.1725 ;
      END
   END din0[118]
   PIN din0[119]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  502.03 1.0375 502.165 1.1725 ;
      END
   END din0[119]
   PIN din0[120]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  504.89 1.0375 505.025 1.1725 ;
      END
   END din0[120]
   PIN din0[121]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  507.75 1.0375 507.885 1.1725 ;
      END
   END din0[121]
   PIN din0[122]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  510.61 1.0375 510.745 1.1725 ;
      END
   END din0[122]
   PIN din0[123]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  513.47 1.0375 513.605 1.1725 ;
      END
   END din0[123]
   PIN din0[124]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  516.33 1.0375 516.465 1.1725 ;
      END
   END din0[124]
   PIN din0[125]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  519.19 1.0375 519.325 1.1725 ;
      END
   END din0[125]
   PIN din0[126]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  522.05 1.0375 522.185 1.1725 ;
      END
   END din0[126]
   PIN din0[127]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  524.91 1.0375 525.045 1.1725 ;
      END
   END din0[127]
   PIN din0[128]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  527.77 1.0375 527.905 1.1725 ;
      END
   END din0[128]
   PIN din0[129]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  530.63 1.0375 530.765 1.1725 ;
      END
   END din0[129]
   PIN din0[130]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  533.49 1.0375 533.625 1.1725 ;
      END
   END din0[130]
   PIN din0[131]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  536.35 1.0375 536.485 1.1725 ;
      END
   END din0[131]
   PIN din0[132]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  539.21 1.0375 539.345 1.1725 ;
      END
   END din0[132]
   PIN din0[133]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  542.07 1.0375 542.205 1.1725 ;
      END
   END din0[133]
   PIN din0[134]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  544.93 1.0375 545.065 1.1725 ;
      END
   END din0[134]
   PIN din0[135]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  547.79 1.0375 547.925 1.1725 ;
      END
   END din0[135]
   PIN din0[136]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  550.65 1.0375 550.785 1.1725 ;
      END
   END din0[136]
   PIN din0[137]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  553.51 1.0375 553.645 1.1725 ;
      END
   END din0[137]
   PIN din0[138]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  556.37 1.0375 556.505 1.1725 ;
      END
   END din0[138]
   PIN din0[139]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  559.23 1.0375 559.365 1.1725 ;
      END
   END din0[139]
   PIN din0[140]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  562.09 1.0375 562.225 1.1725 ;
      END
   END din0[140]
   PIN din0[141]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  564.95 1.0375 565.085 1.1725 ;
      END
   END din0[141]
   PIN din0[142]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  567.81 1.0375 567.945 1.1725 ;
      END
   END din0[142]
   PIN din0[143]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  570.67 1.0375 570.805 1.1725 ;
      END
   END din0[143]
   PIN din0[144]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  573.53 1.0375 573.665 1.1725 ;
      END
   END din0[144]
   PIN din0[145]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  576.39 1.0375 576.525 1.1725 ;
      END
   END din0[145]
   PIN din0[146]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  579.25 1.0375 579.385 1.1725 ;
      END
   END din0[146]
   PIN din0[147]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  582.11 1.0375 582.245 1.1725 ;
      END
   END din0[147]
   PIN din0[148]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  584.97 1.0375 585.105 1.1725 ;
      END
   END din0[148]
   PIN din0[149]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  587.83 1.0375 587.965 1.1725 ;
      END
   END din0[149]
   PIN din0[150]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  590.69 1.0375 590.825 1.1725 ;
      END
   END din0[150]
   PIN din0[151]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  593.55 1.0375 593.685 1.1725 ;
      END
   END din0[151]
   PIN din0[152]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  596.41 1.0375 596.545 1.1725 ;
      END
   END din0[152]
   PIN din0[153]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  599.27 1.0375 599.405 1.1725 ;
      END
   END din0[153]
   PIN din0[154]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  602.13 1.0375 602.265 1.1725 ;
      END
   END din0[154]
   PIN din0[155]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  604.99 1.0375 605.125 1.1725 ;
      END
   END din0[155]
   PIN din0[156]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  607.85 1.0375 607.985 1.1725 ;
      END
   END din0[156]
   PIN din0[157]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  610.71 1.0375 610.845 1.1725 ;
      END
   END din0[157]
   PIN din0[158]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  613.57 1.0375 613.705 1.1725 ;
      END
   END din0[158]
   PIN din0[159]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  616.43 1.0375 616.565 1.1725 ;
      END
   END din0[159]
   PIN din0[160]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  619.29 1.0375 619.425 1.1725 ;
      END
   END din0[160]
   PIN din0[161]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  622.15 1.0375 622.285 1.1725 ;
      END
   END din0[161]
   PIN din0[162]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  625.01 1.0375 625.145 1.1725 ;
      END
   END din0[162]
   PIN din0[163]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  627.87 1.0375 628.005 1.1725 ;
      END
   END din0[163]
   PIN din0[164]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  630.73 1.0375 630.865 1.1725 ;
      END
   END din0[164]
   PIN din0[165]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  633.59 1.0375 633.725 1.1725 ;
      END
   END din0[165]
   PIN din0[166]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  636.45 1.0375 636.585 1.1725 ;
      END
   END din0[166]
   PIN din0[167]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  639.31 1.0375 639.445 1.1725 ;
      END
   END din0[167]
   PIN din0[168]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  642.17 1.0375 642.305 1.1725 ;
      END
   END din0[168]
   PIN din0[169]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  645.03 1.0375 645.165 1.1725 ;
      END
   END din0[169]
   PIN din0[170]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  647.89 1.0375 648.025 1.1725 ;
      END
   END din0[170]
   PIN din0[171]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  650.75 1.0375 650.885 1.1725 ;
      END
   END din0[171]
   PIN din0[172]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  653.61 1.0375 653.745 1.1725 ;
      END
   END din0[172]
   PIN din0[173]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  656.47 1.0375 656.605 1.1725 ;
      END
   END din0[173]
   PIN din0[174]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  659.33 1.0375 659.465 1.1725 ;
      END
   END din0[174]
   PIN din0[175]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  662.19 1.0375 662.325 1.1725 ;
      END
   END din0[175]
   PIN din0[176]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  665.05 1.0375 665.185 1.1725 ;
      END
   END din0[176]
   PIN din0[177]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  667.91 1.0375 668.045 1.1725 ;
      END
   END din0[177]
   PIN din0[178]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  670.77 1.0375 670.905 1.1725 ;
      END
   END din0[178]
   PIN din0[179]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  673.63 1.0375 673.765 1.1725 ;
      END
   END din0[179]
   PIN din0[180]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  676.49 1.0375 676.625 1.1725 ;
      END
   END din0[180]
   PIN din0[181]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  679.35 1.0375 679.485 1.1725 ;
      END
   END din0[181]
   PIN din0[182]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  682.21 1.0375 682.345 1.1725 ;
      END
   END din0[182]
   PIN din0[183]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  685.07 1.0375 685.205 1.1725 ;
      END
   END din0[183]
   PIN din0[184]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  687.93 1.0375 688.065 1.1725 ;
      END
   END din0[184]
   PIN din0[185]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  690.79 1.0375 690.925 1.1725 ;
      END
   END din0[185]
   PIN din0[186]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  693.65 1.0375 693.785 1.1725 ;
      END
   END din0[186]
   PIN din0[187]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  696.51 1.0375 696.645 1.1725 ;
      END
   END din0[187]
   PIN din0[188]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  699.37 1.0375 699.505 1.1725 ;
      END
   END din0[188]
   PIN din0[189]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  702.23 1.0375 702.365 1.1725 ;
      END
   END din0[189]
   PIN din0[190]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  705.09 1.0375 705.225 1.1725 ;
      END
   END din0[190]
   PIN din0[191]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  707.95 1.0375 708.085 1.1725 ;
      END
   END din0[191]
   PIN din0[192]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  710.81 1.0375 710.945 1.1725 ;
      END
   END din0[192]
   PIN din0[193]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  713.67 1.0375 713.805 1.1725 ;
      END
   END din0[193]
   PIN din0[194]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  716.53 1.0375 716.665 1.1725 ;
      END
   END din0[194]
   PIN din0[195]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  719.39 1.0375 719.525 1.1725 ;
      END
   END din0[195]
   PIN din0[196]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  722.25 1.0375 722.385 1.1725 ;
      END
   END din0[196]
   PIN din0[197]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  725.11 1.0375 725.245 1.1725 ;
      END
   END din0[197]
   PIN din0[198]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  727.97 1.0375 728.105 1.1725 ;
      END
   END din0[198]
   PIN din0[199]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  730.83 1.0375 730.965 1.1725 ;
      END
   END din0[199]
   PIN din0[200]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  733.69 1.0375 733.825 1.1725 ;
      END
   END din0[200]
   PIN din0[201]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  736.55 1.0375 736.685 1.1725 ;
      END
   END din0[201]
   PIN din0[202]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  739.41 1.0375 739.545 1.1725 ;
      END
   END din0[202]
   PIN din0[203]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  742.27 1.0375 742.405 1.1725 ;
      END
   END din0[203]
   PIN din0[204]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  745.13 1.0375 745.265 1.1725 ;
      END
   END din0[204]
   PIN din0[205]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  747.99 1.0375 748.125 1.1725 ;
      END
   END din0[205]
   PIN din0[206]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  750.85 1.0375 750.985 1.1725 ;
      END
   END din0[206]
   PIN din0[207]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  753.71 1.0375 753.845 1.1725 ;
      END
   END din0[207]
   PIN din0[208]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  756.57 1.0375 756.705 1.1725 ;
      END
   END din0[208]
   PIN din0[209]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  759.43 1.0375 759.565 1.1725 ;
      END
   END din0[209]
   PIN din0[210]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  762.29 1.0375 762.425 1.1725 ;
      END
   END din0[210]
   PIN din0[211]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  765.15 1.0375 765.285 1.1725 ;
      END
   END din0[211]
   PIN din0[212]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  768.01 1.0375 768.145 1.1725 ;
      END
   END din0[212]
   PIN din0[213]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  770.87 1.0375 771.005 1.1725 ;
      END
   END din0[213]
   PIN din0[214]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  773.73 1.0375 773.865 1.1725 ;
      END
   END din0[214]
   PIN din0[215]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  776.59 1.0375 776.725 1.1725 ;
      END
   END din0[215]
   PIN din0[216]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  779.45 1.0375 779.585 1.1725 ;
      END
   END din0[216]
   PIN din0[217]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  782.31 1.0375 782.445 1.1725 ;
      END
   END din0[217]
   PIN din0[218]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  785.17 1.0375 785.305 1.1725 ;
      END
   END din0[218]
   PIN din0[219]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  788.03 1.0375 788.165 1.1725 ;
      END
   END din0[219]
   PIN din0[220]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  790.89 1.0375 791.025 1.1725 ;
      END
   END din0[220]
   PIN din0[221]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  793.75 1.0375 793.885 1.1725 ;
      END
   END din0[221]
   PIN din0[222]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  796.61 1.0375 796.745 1.1725 ;
      END
   END din0[222]
   PIN din0[223]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  799.47 1.0375 799.605 1.1725 ;
      END
   END din0[223]
   PIN din0[224]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  802.33 1.0375 802.465 1.1725 ;
      END
   END din0[224]
   PIN din0[225]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  805.19 1.0375 805.325 1.1725 ;
      END
   END din0[225]
   PIN din0[226]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  808.05 1.0375 808.185 1.1725 ;
      END
   END din0[226]
   PIN din0[227]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  810.91 1.0375 811.045 1.1725 ;
      END
   END din0[227]
   PIN din0[228]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  813.77 1.0375 813.905 1.1725 ;
      END
   END din0[228]
   PIN din0[229]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  816.63 1.0375 816.765 1.1725 ;
      END
   END din0[229]
   PIN din0[230]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  819.49 1.0375 819.625 1.1725 ;
      END
   END din0[230]
   PIN din0[231]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  822.35 1.0375 822.485 1.1725 ;
      END
   END din0[231]
   PIN din0[232]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  825.21 1.0375 825.345 1.1725 ;
      END
   END din0[232]
   PIN din0[233]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  828.07 1.0375 828.205 1.1725 ;
      END
   END din0[233]
   PIN din0[234]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  830.93 1.0375 831.065 1.1725 ;
      END
   END din0[234]
   PIN din0[235]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  833.79 1.0375 833.925 1.1725 ;
      END
   END din0[235]
   PIN din0[236]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  836.65 1.0375 836.785 1.1725 ;
      END
   END din0[236]
   PIN din0[237]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  839.51 1.0375 839.645 1.1725 ;
      END
   END din0[237]
   PIN din0[238]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  842.37 1.0375 842.505 1.1725 ;
      END
   END din0[238]
   PIN din0[239]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  845.23 1.0375 845.365 1.1725 ;
      END
   END din0[239]
   PIN din0[240]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  848.09 1.0375 848.225 1.1725 ;
      END
   END din0[240]
   PIN din0[241]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  850.95 1.0375 851.085 1.1725 ;
      END
   END din0[241]
   PIN din0[242]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  853.81 1.0375 853.945 1.1725 ;
      END
   END din0[242]
   PIN din0[243]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  856.67 1.0375 856.805 1.1725 ;
      END
   END din0[243]
   PIN din0[244]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  859.53 1.0375 859.665 1.1725 ;
      END
   END din0[244]
   PIN din0[245]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  862.39 1.0375 862.525 1.1725 ;
      END
   END din0[245]
   PIN din0[246]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  865.25 1.0375 865.385 1.1725 ;
      END
   END din0[246]
   PIN din0[247]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  868.11 1.0375 868.245 1.1725 ;
      END
   END din0[247]
   PIN din0[248]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  870.97 1.0375 871.105 1.1725 ;
      END
   END din0[248]
   PIN din0[249]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  873.83 1.0375 873.965 1.1725 ;
      END
   END din0[249]
   PIN din0[250]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  876.69 1.0375 876.825 1.1725 ;
      END
   END din0[250]
   PIN din0[251]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  879.55 1.0375 879.685 1.1725 ;
      END
   END din0[251]
   PIN din0[252]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  882.41 1.0375 882.545 1.1725 ;
      END
   END din0[252]
   PIN din0[253]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  885.27 1.0375 885.405 1.1725 ;
      END
   END din0[253]
   PIN din0[254]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  888.13 1.0375 888.265 1.1725 ;
      END
   END din0[254]
   PIN din0[255]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  890.99 1.0375 891.125 1.1725 ;
      END
   END din0[255]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.45 102.35 64.585 102.485 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.45 105.08 64.585 105.215 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.45 107.29 64.585 107.425 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.45 110.02 64.585 110.155 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.45 112.23 64.585 112.365 ;
      END
   END addr0[4]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 60.36 0.42 60.495 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 63.09 0.42 63.225 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.5275 60.445 6.6625 60.58 ;
      END
   END clk0
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.17 1.0375 70.305 1.1725 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.03 1.0375 73.165 1.1725 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.89 1.0375 76.025 1.1725 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.75 1.0375 78.885 1.1725 ;
      END
   END wmask0[3]
   PIN wmask0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.61 1.0375 81.745 1.1725 ;
      END
   END wmask0[4]
   PIN wmask0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  84.47 1.0375 84.605 1.1725 ;
      END
   END wmask0[5]
   PIN wmask0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  87.33 1.0375 87.465 1.1725 ;
      END
   END wmask0[6]
   PIN wmask0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.19 1.0375 90.325 1.1725 ;
      END
   END wmask0[7]
   PIN wmask0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  93.05 1.0375 93.185 1.1725 ;
      END
   END wmask0[8]
   PIN wmask0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.91 1.0375 96.045 1.1725 ;
      END
   END wmask0[9]
   PIN wmask0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.77 1.0375 98.905 1.1725 ;
      END
   END wmask0[10]
   PIN wmask0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.63 1.0375 101.765 1.1725 ;
      END
   END wmask0[11]
   PIN wmask0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.49 1.0375 104.625 1.1725 ;
      END
   END wmask0[12]
   PIN wmask0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  107.35 1.0375 107.485 1.1725 ;
      END
   END wmask0[13]
   PIN wmask0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  110.21 1.0375 110.345 1.1725 ;
      END
   END wmask0[14]
   PIN wmask0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.07 1.0375 113.205 1.1725 ;
      END
   END wmask0[15]
   PIN wmask0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  115.93 1.0375 116.065 1.1725 ;
      END
   END wmask0[16]
   PIN wmask0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.79 1.0375 118.925 1.1725 ;
      END
   END wmask0[17]
   PIN wmask0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  121.65 1.0375 121.785 1.1725 ;
      END
   END wmask0[18]
   PIN wmask0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  124.51 1.0375 124.645 1.1725 ;
      END
   END wmask0[19]
   PIN wmask0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  127.37 1.0375 127.505 1.1725 ;
      END
   END wmask0[20]
   PIN wmask0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  130.23 1.0375 130.365 1.1725 ;
      END
   END wmask0[21]
   PIN wmask0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  133.09 1.0375 133.225 1.1725 ;
      END
   END wmask0[22]
   PIN wmask0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.95 1.0375 136.085 1.1725 ;
      END
   END wmask0[23]
   PIN wmask0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  138.81 1.0375 138.945 1.1725 ;
      END
   END wmask0[24]
   PIN wmask0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  141.67 1.0375 141.805 1.1725 ;
      END
   END wmask0[25]
   PIN wmask0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  144.53 1.0375 144.665 1.1725 ;
      END
   END wmask0[26]
   PIN wmask0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  147.39 1.0375 147.525 1.1725 ;
      END
   END wmask0[27]
   PIN wmask0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  150.25 1.0375 150.385 1.1725 ;
      END
   END wmask0[28]
   PIN wmask0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  153.11 1.0375 153.245 1.1725 ;
      END
   END wmask0[29]
   PIN wmask0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  155.97 1.0375 156.105 1.1725 ;
      END
   END wmask0[30]
   PIN wmask0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  158.83 1.0375 158.965 1.1725 ;
      END
   END wmask0[31]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.285 71.5025 94.42 71.6375 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.99 71.5025 95.125 71.6375 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.695 71.5025 95.83 71.6375 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.4 71.5025 96.535 71.6375 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.105 71.5025 97.24 71.6375 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.81 71.5025 97.945 71.6375 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.515 71.5025 98.65 71.6375 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.22 71.5025 99.355 71.6375 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.925 71.5025 100.06 71.6375 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.63 71.5025 100.765 71.6375 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.335 71.5025 101.47 71.6375 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  102.04 71.5025 102.175 71.6375 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  102.745 71.5025 102.88 71.6375 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.45 71.5025 103.585 71.6375 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.155 71.5025 104.29 71.6375 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.86 71.5025 104.995 71.6375 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  105.565 71.5025 105.7 71.6375 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.27 71.5025 106.405 71.6375 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.975 71.5025 107.11 71.6375 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  107.68 71.5025 107.815 71.6375 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.385 71.5025 108.52 71.6375 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.09 71.5025 109.225 71.6375 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.795 71.5025 109.93 71.6375 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  110.5 71.5025 110.635 71.6375 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.205 71.5025 111.34 71.6375 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.91 71.5025 112.045 71.6375 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  112.615 71.5025 112.75 71.6375 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.32 71.5025 113.455 71.6375 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.025 71.5025 114.16 71.6375 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.73 71.5025 114.865 71.6375 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  115.435 71.5025 115.57 71.6375 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  116.14 71.5025 116.275 71.6375 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  116.845 71.5025 116.98 71.6375 ;
      END
   END dout0[32]
   PIN dout0[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  117.55 71.5025 117.685 71.6375 ;
      END
   END dout0[33]
   PIN dout0[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.255 71.5025 118.39 71.6375 ;
      END
   END dout0[34]
   PIN dout0[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.96 71.5025 119.095 71.6375 ;
      END
   END dout0[35]
   PIN dout0[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  119.665 71.5025 119.8 71.6375 ;
      END
   END dout0[36]
   PIN dout0[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.37 71.5025 120.505 71.6375 ;
      END
   END dout0[37]
   PIN dout0[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  121.075 71.5025 121.21 71.6375 ;
      END
   END dout0[38]
   PIN dout0[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  121.78 71.5025 121.915 71.6375 ;
      END
   END dout0[39]
   PIN dout0[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  122.485 71.5025 122.62 71.6375 ;
      END
   END dout0[40]
   PIN dout0[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.19 71.5025 123.325 71.6375 ;
      END
   END dout0[41]
   PIN dout0[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.895 71.5025 124.03 71.6375 ;
      END
   END dout0[42]
   PIN dout0[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  124.6 71.5025 124.735 71.6375 ;
      END
   END dout0[43]
   PIN dout0[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  125.305 71.5025 125.44 71.6375 ;
      END
   END dout0[44]
   PIN dout0[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.01 71.5025 126.145 71.6375 ;
      END
   END dout0[45]
   PIN dout0[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.715 71.5025 126.85 71.6375 ;
      END
   END dout0[46]
   PIN dout0[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  127.42 71.5025 127.555 71.6375 ;
      END
   END dout0[47]
   PIN dout0[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  128.125 71.5025 128.26 71.6375 ;
      END
   END dout0[48]
   PIN dout0[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  128.83 71.5025 128.965 71.6375 ;
      END
   END dout0[49]
   PIN dout0[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.535 71.5025 129.67 71.6375 ;
      END
   END dout0[50]
   PIN dout0[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  130.24 71.5025 130.375 71.6375 ;
      END
   END dout0[51]
   PIN dout0[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  130.945 71.5025 131.08 71.6375 ;
      END
   END dout0[52]
   PIN dout0[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.65 71.5025 131.785 71.6375 ;
      END
   END dout0[53]
   PIN dout0[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.355 71.5025 132.49 71.6375 ;
      END
   END dout0[54]
   PIN dout0[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  133.06 71.5025 133.195 71.6375 ;
      END
   END dout0[55]
   PIN dout0[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  133.765 71.5025 133.9 71.6375 ;
      END
   END dout0[56]
   PIN dout0[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.47 71.5025 134.605 71.6375 ;
      END
   END dout0[57]
   PIN dout0[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.175 71.5025 135.31 71.6375 ;
      END
   END dout0[58]
   PIN dout0[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.88 71.5025 136.015 71.6375 ;
      END
   END dout0[59]
   PIN dout0[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  136.585 71.5025 136.72 71.6375 ;
      END
   END dout0[60]
   PIN dout0[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.29 71.5025 137.425 71.6375 ;
      END
   END dout0[61]
   PIN dout0[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.995 71.5025 138.13 71.6375 ;
      END
   END dout0[62]
   PIN dout0[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  138.7 71.5025 138.835 71.6375 ;
      END
   END dout0[63]
   PIN dout0[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  139.405 71.5025 139.54 71.6375 ;
      END
   END dout0[64]
   PIN dout0[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.11 71.5025 140.245 71.6375 ;
      END
   END dout0[65]
   PIN dout0[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.815 71.5025 140.95 71.6375 ;
      END
   END dout0[66]
   PIN dout0[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  141.52 71.5025 141.655 71.6375 ;
      END
   END dout0[67]
   PIN dout0[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  142.225 71.5025 142.36 71.6375 ;
      END
   END dout0[68]
   PIN dout0[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  142.93 71.5025 143.065 71.6375 ;
      END
   END dout0[69]
   PIN dout0[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.635 71.5025 143.77 71.6375 ;
      END
   END dout0[70]
   PIN dout0[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  144.34 71.5025 144.475 71.6375 ;
      END
   END dout0[71]
   PIN dout0[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  145.045 71.5025 145.18 71.6375 ;
      END
   END dout0[72]
   PIN dout0[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  145.75 71.5025 145.885 71.6375 ;
      END
   END dout0[73]
   PIN dout0[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.455 71.5025 146.59 71.6375 ;
      END
   END dout0[74]
   PIN dout0[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  147.16 71.5025 147.295 71.6375 ;
      END
   END dout0[75]
   PIN dout0[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  147.865 71.5025 148.0 71.6375 ;
      END
   END dout0[76]
   PIN dout0[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  148.57 71.5025 148.705 71.6375 ;
      END
   END dout0[77]
   PIN dout0[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.275 71.5025 149.41 71.6375 ;
      END
   END dout0[78]
   PIN dout0[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.98 71.5025 150.115 71.6375 ;
      END
   END dout0[79]
   PIN dout0[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  150.685 71.5025 150.82 71.6375 ;
      END
   END dout0[80]
   PIN dout0[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  151.39 71.5025 151.525 71.6375 ;
      END
   END dout0[81]
   PIN dout0[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.095 71.5025 152.23 71.6375 ;
      END
   END dout0[82]
   PIN dout0[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.8 71.5025 152.935 71.6375 ;
      END
   END dout0[83]
   PIN dout0[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  153.505 71.5025 153.64 71.6375 ;
      END
   END dout0[84]
   PIN dout0[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.21 71.5025 154.345 71.6375 ;
      END
   END dout0[85]
   PIN dout0[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.915 71.5025 155.05 71.6375 ;
      END
   END dout0[86]
   PIN dout0[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  155.62 71.5025 155.755 71.6375 ;
      END
   END dout0[87]
   PIN dout0[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  156.325 71.5025 156.46 71.6375 ;
      END
   END dout0[88]
   PIN dout0[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  157.03 71.5025 157.165 71.6375 ;
      END
   END dout0[89]
   PIN dout0[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  157.735 71.5025 157.87 71.6375 ;
      END
   END dout0[90]
   PIN dout0[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  158.44 71.5025 158.575 71.6375 ;
      END
   END dout0[91]
   PIN dout0[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  159.145 71.5025 159.28 71.6375 ;
      END
   END dout0[92]
   PIN dout0[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  159.85 71.5025 159.985 71.6375 ;
      END
   END dout0[93]
   PIN dout0[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.555 71.5025 160.69 71.6375 ;
      END
   END dout0[94]
   PIN dout0[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  161.26 71.5025 161.395 71.6375 ;
      END
   END dout0[95]
   PIN dout0[96]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  161.965 71.5025 162.1 71.6375 ;
      END
   END dout0[96]
   PIN dout0[97]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  162.67 71.5025 162.805 71.6375 ;
      END
   END dout0[97]
   PIN dout0[98]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.375 71.5025 163.51 71.6375 ;
      END
   END dout0[98]
   PIN dout0[99]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  164.08 71.5025 164.215 71.6375 ;
      END
   END dout0[99]
   PIN dout0[100]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  164.785 71.5025 164.92 71.6375 ;
      END
   END dout0[100]
   PIN dout0[101]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  165.49 71.5025 165.625 71.6375 ;
      END
   END dout0[101]
   PIN dout0[102]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.195 71.5025 166.33 71.6375 ;
      END
   END dout0[102]
   PIN dout0[103]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.9 71.5025 167.035 71.6375 ;
      END
   END dout0[103]
   PIN dout0[104]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  167.605 71.5025 167.74 71.6375 ;
      END
   END dout0[104]
   PIN dout0[105]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  168.31 71.5025 168.445 71.6375 ;
      END
   END dout0[105]
   PIN dout0[106]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.015 71.5025 169.15 71.6375 ;
      END
   END dout0[106]
   PIN dout0[107]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.72 71.5025 169.855 71.6375 ;
      END
   END dout0[107]
   PIN dout0[108]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  170.425 71.5025 170.56 71.6375 ;
      END
   END dout0[108]
   PIN dout0[109]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  171.13 71.5025 171.265 71.6375 ;
      END
   END dout0[109]
   PIN dout0[110]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  171.835 71.5025 171.97 71.6375 ;
      END
   END dout0[110]
   PIN dout0[111]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.54 71.5025 172.675 71.6375 ;
      END
   END dout0[111]
   PIN dout0[112]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  173.245 71.5025 173.38 71.6375 ;
      END
   END dout0[112]
   PIN dout0[113]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  173.95 71.5025 174.085 71.6375 ;
      END
   END dout0[113]
   PIN dout0[114]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.655 71.5025 174.79 71.6375 ;
      END
   END dout0[114]
   PIN dout0[115]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  175.36 71.5025 175.495 71.6375 ;
      END
   END dout0[115]
   PIN dout0[116]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  176.065 71.5025 176.2 71.6375 ;
      END
   END dout0[116]
   PIN dout0[117]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  176.77 71.5025 176.905 71.6375 ;
      END
   END dout0[117]
   PIN dout0[118]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.475 71.5025 177.61 71.6375 ;
      END
   END dout0[118]
   PIN dout0[119]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.18 71.5025 178.315 71.6375 ;
      END
   END dout0[119]
   PIN dout0[120]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.885 71.5025 179.02 71.6375 ;
      END
   END dout0[120]
   PIN dout0[121]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.59 71.5025 179.725 71.6375 ;
      END
   END dout0[121]
   PIN dout0[122]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.295 71.5025 180.43 71.6375 ;
      END
   END dout0[122]
   PIN dout0[123]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  181.0 71.5025 181.135 71.6375 ;
      END
   END dout0[123]
   PIN dout0[124]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  181.705 71.5025 181.84 71.6375 ;
      END
   END dout0[124]
   PIN dout0[125]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  182.41 71.5025 182.545 71.6375 ;
      END
   END dout0[125]
   PIN dout0[126]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.115 71.5025 183.25 71.6375 ;
      END
   END dout0[126]
   PIN dout0[127]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.82 71.5025 183.955 71.6375 ;
      END
   END dout0[127]
   PIN dout0[128]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  184.525 71.5025 184.66 71.6375 ;
      END
   END dout0[128]
   PIN dout0[129]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.23 71.5025 185.365 71.6375 ;
      END
   END dout0[129]
   PIN dout0[130]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.935 71.5025 186.07 71.6375 ;
      END
   END dout0[130]
   PIN dout0[131]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.64 71.5025 186.775 71.6375 ;
      END
   END dout0[131]
   PIN dout0[132]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  187.345 71.5025 187.48 71.6375 ;
      END
   END dout0[132]
   PIN dout0[133]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  188.05 71.5025 188.185 71.6375 ;
      END
   END dout0[133]
   PIN dout0[134]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  188.755 71.5025 188.89 71.6375 ;
      END
   END dout0[134]
   PIN dout0[135]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.46 71.5025 189.595 71.6375 ;
      END
   END dout0[135]
   PIN dout0[136]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  190.165 71.5025 190.3 71.6375 ;
      END
   END dout0[136]
   PIN dout0[137]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  190.87 71.5025 191.005 71.6375 ;
      END
   END dout0[137]
   PIN dout0[138]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  191.575 71.5025 191.71 71.6375 ;
      END
   END dout0[138]
   PIN dout0[139]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.28 71.5025 192.415 71.6375 ;
      END
   END dout0[139]
   PIN dout0[140]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.985 71.5025 193.12 71.6375 ;
      END
   END dout0[140]
   PIN dout0[141]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  193.69 71.5025 193.825 71.6375 ;
      END
   END dout0[141]
   PIN dout0[142]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  194.395 71.5025 194.53 71.6375 ;
      END
   END dout0[142]
   PIN dout0[143]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  195.1 71.5025 195.235 71.6375 ;
      END
   END dout0[143]
   PIN dout0[144]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  195.805 71.5025 195.94 71.6375 ;
      END
   END dout0[144]
   PIN dout0[145]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  196.51 71.5025 196.645 71.6375 ;
      END
   END dout0[145]
   PIN dout0[146]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  197.215 71.5025 197.35 71.6375 ;
      END
   END dout0[146]
   PIN dout0[147]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  197.92 71.5025 198.055 71.6375 ;
      END
   END dout0[147]
   PIN dout0[148]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  198.625 71.5025 198.76 71.6375 ;
      END
   END dout0[148]
   PIN dout0[149]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  199.33 71.5025 199.465 71.6375 ;
      END
   END dout0[149]
   PIN dout0[150]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  200.035 71.5025 200.17 71.6375 ;
      END
   END dout0[150]
   PIN dout0[151]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  200.74 71.5025 200.875 71.6375 ;
      END
   END dout0[151]
   PIN dout0[152]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  201.445 71.5025 201.58 71.6375 ;
      END
   END dout0[152]
   PIN dout0[153]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  202.15 71.5025 202.285 71.6375 ;
      END
   END dout0[153]
   PIN dout0[154]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  202.855 71.5025 202.99 71.6375 ;
      END
   END dout0[154]
   PIN dout0[155]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  203.56 71.5025 203.695 71.6375 ;
      END
   END dout0[155]
   PIN dout0[156]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  204.265 71.5025 204.4 71.6375 ;
      END
   END dout0[156]
   PIN dout0[157]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  204.97 71.5025 205.105 71.6375 ;
      END
   END dout0[157]
   PIN dout0[158]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  205.675 71.5025 205.81 71.6375 ;
      END
   END dout0[158]
   PIN dout0[159]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  206.38 71.5025 206.515 71.6375 ;
      END
   END dout0[159]
   PIN dout0[160]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  207.085 71.5025 207.22 71.6375 ;
      END
   END dout0[160]
   PIN dout0[161]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  207.79 71.5025 207.925 71.6375 ;
      END
   END dout0[161]
   PIN dout0[162]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  208.495 71.5025 208.63 71.6375 ;
      END
   END dout0[162]
   PIN dout0[163]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  209.2 71.5025 209.335 71.6375 ;
      END
   END dout0[163]
   PIN dout0[164]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  209.905 71.5025 210.04 71.6375 ;
      END
   END dout0[164]
   PIN dout0[165]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  210.61 71.5025 210.745 71.6375 ;
      END
   END dout0[165]
   PIN dout0[166]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  211.315 71.5025 211.45 71.6375 ;
      END
   END dout0[166]
   PIN dout0[167]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.02 71.5025 212.155 71.6375 ;
      END
   END dout0[167]
   PIN dout0[168]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.725 71.5025 212.86 71.6375 ;
      END
   END dout0[168]
   PIN dout0[169]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  213.43 71.5025 213.565 71.6375 ;
      END
   END dout0[169]
   PIN dout0[170]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  214.135 71.5025 214.27 71.6375 ;
      END
   END dout0[170]
   PIN dout0[171]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  214.84 71.5025 214.975 71.6375 ;
      END
   END dout0[171]
   PIN dout0[172]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  215.545 71.5025 215.68 71.6375 ;
      END
   END dout0[172]
   PIN dout0[173]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  216.25 71.5025 216.385 71.6375 ;
      END
   END dout0[173]
   PIN dout0[174]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  216.955 71.5025 217.09 71.6375 ;
      END
   END dout0[174]
   PIN dout0[175]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  217.66 71.5025 217.795 71.6375 ;
      END
   END dout0[175]
   PIN dout0[176]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  218.365 71.5025 218.5 71.6375 ;
      END
   END dout0[176]
   PIN dout0[177]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  219.07 71.5025 219.205 71.6375 ;
      END
   END dout0[177]
   PIN dout0[178]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  219.775 71.5025 219.91 71.6375 ;
      END
   END dout0[178]
   PIN dout0[179]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  220.48 71.5025 220.615 71.6375 ;
      END
   END dout0[179]
   PIN dout0[180]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  221.185 71.5025 221.32 71.6375 ;
      END
   END dout0[180]
   PIN dout0[181]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  221.89 71.5025 222.025 71.6375 ;
      END
   END dout0[181]
   PIN dout0[182]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  222.595 71.5025 222.73 71.6375 ;
      END
   END dout0[182]
   PIN dout0[183]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  223.3 71.5025 223.435 71.6375 ;
      END
   END dout0[183]
   PIN dout0[184]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  224.005 71.5025 224.14 71.6375 ;
      END
   END dout0[184]
   PIN dout0[185]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  224.71 71.5025 224.845 71.6375 ;
      END
   END dout0[185]
   PIN dout0[186]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  225.415 71.5025 225.55 71.6375 ;
      END
   END dout0[186]
   PIN dout0[187]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  226.12 71.5025 226.255 71.6375 ;
      END
   END dout0[187]
   PIN dout0[188]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  226.825 71.5025 226.96 71.6375 ;
      END
   END dout0[188]
   PIN dout0[189]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  227.53 71.5025 227.665 71.6375 ;
      END
   END dout0[189]
   PIN dout0[190]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  228.235 71.5025 228.37 71.6375 ;
      END
   END dout0[190]
   PIN dout0[191]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  228.94 71.5025 229.075 71.6375 ;
      END
   END dout0[191]
   PIN dout0[192]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  229.645 71.5025 229.78 71.6375 ;
      END
   END dout0[192]
   PIN dout0[193]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  230.35 71.5025 230.485 71.6375 ;
      END
   END dout0[193]
   PIN dout0[194]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  231.055 71.5025 231.19 71.6375 ;
      END
   END dout0[194]
   PIN dout0[195]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  231.76 71.5025 231.895 71.6375 ;
      END
   END dout0[195]
   PIN dout0[196]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  232.465 71.5025 232.6 71.6375 ;
      END
   END dout0[196]
   PIN dout0[197]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  233.17 71.5025 233.305 71.6375 ;
      END
   END dout0[197]
   PIN dout0[198]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  233.875 71.5025 234.01 71.6375 ;
      END
   END dout0[198]
   PIN dout0[199]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  234.58 71.5025 234.715 71.6375 ;
      END
   END dout0[199]
   PIN dout0[200]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  235.285 71.5025 235.42 71.6375 ;
      END
   END dout0[200]
   PIN dout0[201]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  235.99 71.5025 236.125 71.6375 ;
      END
   END dout0[201]
   PIN dout0[202]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  236.695 71.5025 236.83 71.6375 ;
      END
   END dout0[202]
   PIN dout0[203]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  237.4 71.5025 237.535 71.6375 ;
      END
   END dout0[203]
   PIN dout0[204]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  238.105 71.5025 238.24 71.6375 ;
      END
   END dout0[204]
   PIN dout0[205]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  238.81 71.5025 238.945 71.6375 ;
      END
   END dout0[205]
   PIN dout0[206]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  239.515 71.5025 239.65 71.6375 ;
      END
   END dout0[206]
   PIN dout0[207]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  240.22 71.5025 240.355 71.6375 ;
      END
   END dout0[207]
   PIN dout0[208]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  240.925 71.5025 241.06 71.6375 ;
      END
   END dout0[208]
   PIN dout0[209]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  241.63 71.5025 241.765 71.6375 ;
      END
   END dout0[209]
   PIN dout0[210]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  242.335 71.5025 242.47 71.6375 ;
      END
   END dout0[210]
   PIN dout0[211]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  243.04 71.5025 243.175 71.6375 ;
      END
   END dout0[211]
   PIN dout0[212]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  243.745 71.5025 243.88 71.6375 ;
      END
   END dout0[212]
   PIN dout0[213]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  244.45 71.5025 244.585 71.6375 ;
      END
   END dout0[213]
   PIN dout0[214]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  245.155 71.5025 245.29 71.6375 ;
      END
   END dout0[214]
   PIN dout0[215]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  245.86 71.5025 245.995 71.6375 ;
      END
   END dout0[215]
   PIN dout0[216]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  246.565 71.5025 246.7 71.6375 ;
      END
   END dout0[216]
   PIN dout0[217]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  247.27 71.5025 247.405 71.6375 ;
      END
   END dout0[217]
   PIN dout0[218]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  247.975 71.5025 248.11 71.6375 ;
      END
   END dout0[218]
   PIN dout0[219]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  248.68 71.5025 248.815 71.6375 ;
      END
   END dout0[219]
   PIN dout0[220]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  249.385 71.5025 249.52 71.6375 ;
      END
   END dout0[220]
   PIN dout0[221]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  250.09 71.5025 250.225 71.6375 ;
      END
   END dout0[221]
   PIN dout0[222]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  250.795 71.5025 250.93 71.6375 ;
      END
   END dout0[222]
   PIN dout0[223]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  251.5 71.5025 251.635 71.6375 ;
      END
   END dout0[223]
   PIN dout0[224]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  252.205 71.5025 252.34 71.6375 ;
      END
   END dout0[224]
   PIN dout0[225]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  252.91 71.5025 253.045 71.6375 ;
      END
   END dout0[225]
   PIN dout0[226]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  253.615 71.5025 253.75 71.6375 ;
      END
   END dout0[226]
   PIN dout0[227]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  254.32 71.5025 254.455 71.6375 ;
      END
   END dout0[227]
   PIN dout0[228]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  255.025 71.5025 255.16 71.6375 ;
      END
   END dout0[228]
   PIN dout0[229]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  255.73 71.5025 255.865 71.6375 ;
      END
   END dout0[229]
   PIN dout0[230]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  256.435 71.5025 256.57 71.6375 ;
      END
   END dout0[230]
   PIN dout0[231]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  257.14 71.5025 257.275 71.6375 ;
      END
   END dout0[231]
   PIN dout0[232]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  257.845 71.5025 257.98 71.6375 ;
      END
   END dout0[232]
   PIN dout0[233]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  258.55 71.5025 258.685 71.6375 ;
      END
   END dout0[233]
   PIN dout0[234]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  259.255 71.5025 259.39 71.6375 ;
      END
   END dout0[234]
   PIN dout0[235]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  259.96 71.5025 260.095 71.6375 ;
      END
   END dout0[235]
   PIN dout0[236]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  260.665 71.5025 260.8 71.6375 ;
      END
   END dout0[236]
   PIN dout0[237]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  261.37 71.5025 261.505 71.6375 ;
      END
   END dout0[237]
   PIN dout0[238]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  262.075 71.5025 262.21 71.6375 ;
      END
   END dout0[238]
   PIN dout0[239]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  262.78 71.5025 262.915 71.6375 ;
      END
   END dout0[239]
   PIN dout0[240]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  263.485 71.5025 263.62 71.6375 ;
      END
   END dout0[240]
   PIN dout0[241]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  264.19 71.5025 264.325 71.6375 ;
      END
   END dout0[241]
   PIN dout0[242]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  264.895 71.5025 265.03 71.6375 ;
      END
   END dout0[242]
   PIN dout0[243]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  265.6 71.5025 265.735 71.6375 ;
      END
   END dout0[243]
   PIN dout0[244]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  266.305 71.5025 266.44 71.6375 ;
      END
   END dout0[244]
   PIN dout0[245]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  267.01 71.5025 267.145 71.6375 ;
      END
   END dout0[245]
   PIN dout0[246]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  267.715 71.5025 267.85 71.6375 ;
      END
   END dout0[246]
   PIN dout0[247]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  268.42 71.5025 268.555 71.6375 ;
      END
   END dout0[247]
   PIN dout0[248]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  269.125 71.5025 269.26 71.6375 ;
      END
   END dout0[248]
   PIN dout0[249]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  269.83 71.5025 269.965 71.6375 ;
      END
   END dout0[249]
   PIN dout0[250]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  270.535 71.5025 270.67 71.6375 ;
      END
   END dout0[250]
   PIN dout0[251]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  271.24 71.5025 271.375 71.6375 ;
      END
   END dout0[251]
   PIN dout0[252]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  271.945 71.5025 272.08 71.6375 ;
      END
   END dout0[252]
   PIN dout0[253]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  272.65 71.5025 272.785 71.6375 ;
      END
   END dout0[253]
   PIN dout0[254]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  273.355 71.5025 273.49 71.6375 ;
      END
   END dout0[254]
   PIN dout0[255]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  274.06 71.5025 274.195 71.6375 ;
      END
   END dout0[255]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 893.495 127.305 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 893.495 127.305 ;
   LAYER  metal3 ;
      RECT  0.14 0.14 161.55 0.8975 ;
      RECT  161.55 0.14 161.965 0.8975 ;
      RECT  161.965 0.14 893.495 0.8975 ;
      RECT  161.965 0.8975 164.41 1.3125 ;
      RECT  164.825 0.8975 167.27 1.3125 ;
      RECT  167.685 0.8975 170.13 1.3125 ;
      RECT  170.545 0.8975 172.99 1.3125 ;
      RECT  173.405 0.8975 175.85 1.3125 ;
      RECT  176.265 0.8975 178.71 1.3125 ;
      RECT  179.125 0.8975 181.57 1.3125 ;
      RECT  181.985 0.8975 184.43 1.3125 ;
      RECT  184.845 0.8975 187.29 1.3125 ;
      RECT  187.705 0.8975 190.15 1.3125 ;
      RECT  190.565 0.8975 193.01 1.3125 ;
      RECT  193.425 0.8975 195.87 1.3125 ;
      RECT  196.285 0.8975 198.73 1.3125 ;
      RECT  199.145 0.8975 201.59 1.3125 ;
      RECT  202.005 0.8975 204.45 1.3125 ;
      RECT  204.865 0.8975 207.31 1.3125 ;
      RECT  207.725 0.8975 210.17 1.3125 ;
      RECT  210.585 0.8975 213.03 1.3125 ;
      RECT  213.445 0.8975 215.89 1.3125 ;
      RECT  216.305 0.8975 218.75 1.3125 ;
      RECT  219.165 0.8975 221.61 1.3125 ;
      RECT  222.025 0.8975 224.47 1.3125 ;
      RECT  224.885 0.8975 227.33 1.3125 ;
      RECT  227.745 0.8975 230.19 1.3125 ;
      RECT  230.605 0.8975 233.05 1.3125 ;
      RECT  233.465 0.8975 235.91 1.3125 ;
      RECT  236.325 0.8975 238.77 1.3125 ;
      RECT  239.185 0.8975 241.63 1.3125 ;
      RECT  242.045 0.8975 244.49 1.3125 ;
      RECT  244.905 0.8975 247.35 1.3125 ;
      RECT  247.765 0.8975 250.21 1.3125 ;
      RECT  250.625 0.8975 253.07 1.3125 ;
      RECT  253.485 0.8975 255.93 1.3125 ;
      RECT  256.345 0.8975 258.79 1.3125 ;
      RECT  259.205 0.8975 261.65 1.3125 ;
      RECT  262.065 0.8975 264.51 1.3125 ;
      RECT  264.925 0.8975 267.37 1.3125 ;
      RECT  267.785 0.8975 270.23 1.3125 ;
      RECT  270.645 0.8975 273.09 1.3125 ;
      RECT  273.505 0.8975 275.95 1.3125 ;
      RECT  276.365 0.8975 278.81 1.3125 ;
      RECT  279.225 0.8975 281.67 1.3125 ;
      RECT  282.085 0.8975 284.53 1.3125 ;
      RECT  284.945 0.8975 287.39 1.3125 ;
      RECT  287.805 0.8975 290.25 1.3125 ;
      RECT  290.665 0.8975 293.11 1.3125 ;
      RECT  293.525 0.8975 295.97 1.3125 ;
      RECT  296.385 0.8975 298.83 1.3125 ;
      RECT  299.245 0.8975 301.69 1.3125 ;
      RECT  302.105 0.8975 304.55 1.3125 ;
      RECT  304.965 0.8975 307.41 1.3125 ;
      RECT  307.825 0.8975 310.27 1.3125 ;
      RECT  310.685 0.8975 313.13 1.3125 ;
      RECT  313.545 0.8975 315.99 1.3125 ;
      RECT  316.405 0.8975 318.85 1.3125 ;
      RECT  319.265 0.8975 321.71 1.3125 ;
      RECT  322.125 0.8975 324.57 1.3125 ;
      RECT  324.985 0.8975 327.43 1.3125 ;
      RECT  327.845 0.8975 330.29 1.3125 ;
      RECT  330.705 0.8975 333.15 1.3125 ;
      RECT  333.565 0.8975 336.01 1.3125 ;
      RECT  336.425 0.8975 338.87 1.3125 ;
      RECT  339.285 0.8975 341.73 1.3125 ;
      RECT  342.145 0.8975 344.59 1.3125 ;
      RECT  345.005 0.8975 347.45 1.3125 ;
      RECT  347.865 0.8975 350.31 1.3125 ;
      RECT  350.725 0.8975 353.17 1.3125 ;
      RECT  353.585 0.8975 356.03 1.3125 ;
      RECT  356.445 0.8975 358.89 1.3125 ;
      RECT  359.305 0.8975 361.75 1.3125 ;
      RECT  362.165 0.8975 364.61 1.3125 ;
      RECT  365.025 0.8975 367.47 1.3125 ;
      RECT  367.885 0.8975 370.33 1.3125 ;
      RECT  370.745 0.8975 373.19 1.3125 ;
      RECT  373.605 0.8975 376.05 1.3125 ;
      RECT  376.465 0.8975 378.91 1.3125 ;
      RECT  379.325 0.8975 381.77 1.3125 ;
      RECT  382.185 0.8975 384.63 1.3125 ;
      RECT  385.045 0.8975 387.49 1.3125 ;
      RECT  387.905 0.8975 390.35 1.3125 ;
      RECT  390.765 0.8975 393.21 1.3125 ;
      RECT  393.625 0.8975 396.07 1.3125 ;
      RECT  396.485 0.8975 398.93 1.3125 ;
      RECT  399.345 0.8975 401.79 1.3125 ;
      RECT  402.205 0.8975 404.65 1.3125 ;
      RECT  405.065 0.8975 407.51 1.3125 ;
      RECT  407.925 0.8975 410.37 1.3125 ;
      RECT  410.785 0.8975 413.23 1.3125 ;
      RECT  413.645 0.8975 416.09 1.3125 ;
      RECT  416.505 0.8975 418.95 1.3125 ;
      RECT  419.365 0.8975 421.81 1.3125 ;
      RECT  422.225 0.8975 424.67 1.3125 ;
      RECT  425.085 0.8975 427.53 1.3125 ;
      RECT  427.945 0.8975 430.39 1.3125 ;
      RECT  430.805 0.8975 433.25 1.3125 ;
      RECT  433.665 0.8975 436.11 1.3125 ;
      RECT  436.525 0.8975 438.97 1.3125 ;
      RECT  439.385 0.8975 441.83 1.3125 ;
      RECT  442.245 0.8975 444.69 1.3125 ;
      RECT  445.105 0.8975 447.55 1.3125 ;
      RECT  447.965 0.8975 450.41 1.3125 ;
      RECT  450.825 0.8975 453.27 1.3125 ;
      RECT  453.685 0.8975 456.13 1.3125 ;
      RECT  456.545 0.8975 458.99 1.3125 ;
      RECT  459.405 0.8975 461.85 1.3125 ;
      RECT  462.265 0.8975 464.71 1.3125 ;
      RECT  465.125 0.8975 467.57 1.3125 ;
      RECT  467.985 0.8975 470.43 1.3125 ;
      RECT  470.845 0.8975 473.29 1.3125 ;
      RECT  473.705 0.8975 476.15 1.3125 ;
      RECT  476.565 0.8975 479.01 1.3125 ;
      RECT  479.425 0.8975 481.87 1.3125 ;
      RECT  482.285 0.8975 484.73 1.3125 ;
      RECT  485.145 0.8975 487.59 1.3125 ;
      RECT  488.005 0.8975 490.45 1.3125 ;
      RECT  490.865 0.8975 493.31 1.3125 ;
      RECT  493.725 0.8975 496.17 1.3125 ;
      RECT  496.585 0.8975 499.03 1.3125 ;
      RECT  499.445 0.8975 501.89 1.3125 ;
      RECT  502.305 0.8975 504.75 1.3125 ;
      RECT  505.165 0.8975 507.61 1.3125 ;
      RECT  508.025 0.8975 510.47 1.3125 ;
      RECT  510.885 0.8975 513.33 1.3125 ;
      RECT  513.745 0.8975 516.19 1.3125 ;
      RECT  516.605 0.8975 519.05 1.3125 ;
      RECT  519.465 0.8975 521.91 1.3125 ;
      RECT  522.325 0.8975 524.77 1.3125 ;
      RECT  525.185 0.8975 527.63 1.3125 ;
      RECT  528.045 0.8975 530.49 1.3125 ;
      RECT  530.905 0.8975 533.35 1.3125 ;
      RECT  533.765 0.8975 536.21 1.3125 ;
      RECT  536.625 0.8975 539.07 1.3125 ;
      RECT  539.485 0.8975 541.93 1.3125 ;
      RECT  542.345 0.8975 544.79 1.3125 ;
      RECT  545.205 0.8975 547.65 1.3125 ;
      RECT  548.065 0.8975 550.51 1.3125 ;
      RECT  550.925 0.8975 553.37 1.3125 ;
      RECT  553.785 0.8975 556.23 1.3125 ;
      RECT  556.645 0.8975 559.09 1.3125 ;
      RECT  559.505 0.8975 561.95 1.3125 ;
      RECT  562.365 0.8975 564.81 1.3125 ;
      RECT  565.225 0.8975 567.67 1.3125 ;
      RECT  568.085 0.8975 570.53 1.3125 ;
      RECT  570.945 0.8975 573.39 1.3125 ;
      RECT  573.805 0.8975 576.25 1.3125 ;
      RECT  576.665 0.8975 579.11 1.3125 ;
      RECT  579.525 0.8975 581.97 1.3125 ;
      RECT  582.385 0.8975 584.83 1.3125 ;
      RECT  585.245 0.8975 587.69 1.3125 ;
      RECT  588.105 0.8975 590.55 1.3125 ;
      RECT  590.965 0.8975 593.41 1.3125 ;
      RECT  593.825 0.8975 596.27 1.3125 ;
      RECT  596.685 0.8975 599.13 1.3125 ;
      RECT  599.545 0.8975 601.99 1.3125 ;
      RECT  602.405 0.8975 604.85 1.3125 ;
      RECT  605.265 0.8975 607.71 1.3125 ;
      RECT  608.125 0.8975 610.57 1.3125 ;
      RECT  610.985 0.8975 613.43 1.3125 ;
      RECT  613.845 0.8975 616.29 1.3125 ;
      RECT  616.705 0.8975 619.15 1.3125 ;
      RECT  619.565 0.8975 622.01 1.3125 ;
      RECT  622.425 0.8975 624.87 1.3125 ;
      RECT  625.285 0.8975 627.73 1.3125 ;
      RECT  628.145 0.8975 630.59 1.3125 ;
      RECT  631.005 0.8975 633.45 1.3125 ;
      RECT  633.865 0.8975 636.31 1.3125 ;
      RECT  636.725 0.8975 639.17 1.3125 ;
      RECT  639.585 0.8975 642.03 1.3125 ;
      RECT  642.445 0.8975 644.89 1.3125 ;
      RECT  645.305 0.8975 647.75 1.3125 ;
      RECT  648.165 0.8975 650.61 1.3125 ;
      RECT  651.025 0.8975 653.47 1.3125 ;
      RECT  653.885 0.8975 656.33 1.3125 ;
      RECT  656.745 0.8975 659.19 1.3125 ;
      RECT  659.605 0.8975 662.05 1.3125 ;
      RECT  662.465 0.8975 664.91 1.3125 ;
      RECT  665.325 0.8975 667.77 1.3125 ;
      RECT  668.185 0.8975 670.63 1.3125 ;
      RECT  671.045 0.8975 673.49 1.3125 ;
      RECT  673.905 0.8975 676.35 1.3125 ;
      RECT  676.765 0.8975 679.21 1.3125 ;
      RECT  679.625 0.8975 682.07 1.3125 ;
      RECT  682.485 0.8975 684.93 1.3125 ;
      RECT  685.345 0.8975 687.79 1.3125 ;
      RECT  688.205 0.8975 690.65 1.3125 ;
      RECT  691.065 0.8975 693.51 1.3125 ;
      RECT  693.925 0.8975 696.37 1.3125 ;
      RECT  696.785 0.8975 699.23 1.3125 ;
      RECT  699.645 0.8975 702.09 1.3125 ;
      RECT  702.505 0.8975 704.95 1.3125 ;
      RECT  705.365 0.8975 707.81 1.3125 ;
      RECT  708.225 0.8975 710.67 1.3125 ;
      RECT  711.085 0.8975 713.53 1.3125 ;
      RECT  713.945 0.8975 716.39 1.3125 ;
      RECT  716.805 0.8975 719.25 1.3125 ;
      RECT  719.665 0.8975 722.11 1.3125 ;
      RECT  722.525 0.8975 724.97 1.3125 ;
      RECT  725.385 0.8975 727.83 1.3125 ;
      RECT  728.245 0.8975 730.69 1.3125 ;
      RECT  731.105 0.8975 733.55 1.3125 ;
      RECT  733.965 0.8975 736.41 1.3125 ;
      RECT  736.825 0.8975 739.27 1.3125 ;
      RECT  739.685 0.8975 742.13 1.3125 ;
      RECT  742.545 0.8975 744.99 1.3125 ;
      RECT  745.405 0.8975 747.85 1.3125 ;
      RECT  748.265 0.8975 750.71 1.3125 ;
      RECT  751.125 0.8975 753.57 1.3125 ;
      RECT  753.985 0.8975 756.43 1.3125 ;
      RECT  756.845 0.8975 759.29 1.3125 ;
      RECT  759.705 0.8975 762.15 1.3125 ;
      RECT  762.565 0.8975 765.01 1.3125 ;
      RECT  765.425 0.8975 767.87 1.3125 ;
      RECT  768.285 0.8975 770.73 1.3125 ;
      RECT  771.145 0.8975 773.59 1.3125 ;
      RECT  774.005 0.8975 776.45 1.3125 ;
      RECT  776.865 0.8975 779.31 1.3125 ;
      RECT  779.725 0.8975 782.17 1.3125 ;
      RECT  782.585 0.8975 785.03 1.3125 ;
      RECT  785.445 0.8975 787.89 1.3125 ;
      RECT  788.305 0.8975 790.75 1.3125 ;
      RECT  791.165 0.8975 793.61 1.3125 ;
      RECT  794.025 0.8975 796.47 1.3125 ;
      RECT  796.885 0.8975 799.33 1.3125 ;
      RECT  799.745 0.8975 802.19 1.3125 ;
      RECT  802.605 0.8975 805.05 1.3125 ;
      RECT  805.465 0.8975 807.91 1.3125 ;
      RECT  808.325 0.8975 810.77 1.3125 ;
      RECT  811.185 0.8975 813.63 1.3125 ;
      RECT  814.045 0.8975 816.49 1.3125 ;
      RECT  816.905 0.8975 819.35 1.3125 ;
      RECT  819.765 0.8975 822.21 1.3125 ;
      RECT  822.625 0.8975 825.07 1.3125 ;
      RECT  825.485 0.8975 827.93 1.3125 ;
      RECT  828.345 0.8975 830.79 1.3125 ;
      RECT  831.205 0.8975 833.65 1.3125 ;
      RECT  834.065 0.8975 836.51 1.3125 ;
      RECT  836.925 0.8975 839.37 1.3125 ;
      RECT  839.785 0.8975 842.23 1.3125 ;
      RECT  842.645 0.8975 845.09 1.3125 ;
      RECT  845.505 0.8975 847.95 1.3125 ;
      RECT  848.365 0.8975 850.81 1.3125 ;
      RECT  851.225 0.8975 853.67 1.3125 ;
      RECT  854.085 0.8975 856.53 1.3125 ;
      RECT  856.945 0.8975 859.39 1.3125 ;
      RECT  859.805 0.8975 862.25 1.3125 ;
      RECT  862.665 0.8975 865.11 1.3125 ;
      RECT  865.525 0.8975 867.97 1.3125 ;
      RECT  868.385 0.8975 870.83 1.3125 ;
      RECT  871.245 0.8975 873.69 1.3125 ;
      RECT  874.105 0.8975 876.55 1.3125 ;
      RECT  876.965 0.8975 879.41 1.3125 ;
      RECT  879.825 0.8975 882.27 1.3125 ;
      RECT  882.685 0.8975 885.13 1.3125 ;
      RECT  885.545 0.8975 887.99 1.3125 ;
      RECT  888.405 0.8975 890.85 1.3125 ;
      RECT  891.265 0.8975 893.495 1.3125 ;
      RECT  0.14 102.21 64.31 102.625 ;
      RECT  0.14 102.625 64.31 127.305 ;
      RECT  64.31 1.3125 64.725 102.21 ;
      RECT  64.725 102.21 161.55 102.625 ;
      RECT  64.725 102.625 161.55 127.305 ;
      RECT  64.31 102.625 64.725 104.94 ;
      RECT  64.31 105.355 64.725 107.15 ;
      RECT  64.31 107.565 64.725 109.88 ;
      RECT  64.31 110.295 64.725 112.09 ;
      RECT  64.31 112.505 64.725 127.305 ;
      RECT  0.14 1.3125 0.145 60.22 ;
      RECT  0.14 60.22 0.145 60.635 ;
      RECT  0.14 60.635 0.145 102.21 ;
      RECT  0.145 1.3125 0.56 60.22 ;
      RECT  0.56 1.3125 64.31 60.22 ;
      RECT  0.145 60.635 0.56 62.95 ;
      RECT  0.145 63.365 0.56 102.21 ;
      RECT  0.56 60.22 6.3875 60.305 ;
      RECT  0.56 60.305 6.3875 60.635 ;
      RECT  6.3875 60.22 6.8025 60.305 ;
      RECT  6.8025 60.22 64.31 60.305 ;
      RECT  6.8025 60.305 64.31 60.635 ;
      RECT  0.56 60.635 6.3875 60.72 ;
      RECT  0.56 60.72 6.3875 102.21 ;
      RECT  6.3875 60.72 6.8025 102.21 ;
      RECT  6.8025 60.635 64.31 60.72 ;
      RECT  6.8025 60.72 64.31 102.21 ;
      RECT  0.14 0.8975 70.03 1.3125 ;
      RECT  70.445 0.8975 72.89 1.3125 ;
      RECT  73.305 0.8975 75.75 1.3125 ;
      RECT  76.165 0.8975 78.61 1.3125 ;
      RECT  79.025 0.8975 81.47 1.3125 ;
      RECT  81.885 0.8975 84.33 1.3125 ;
      RECT  84.745 0.8975 87.19 1.3125 ;
      RECT  87.605 0.8975 90.05 1.3125 ;
      RECT  90.465 0.8975 92.91 1.3125 ;
      RECT  93.325 0.8975 95.77 1.3125 ;
      RECT  96.185 0.8975 98.63 1.3125 ;
      RECT  99.045 0.8975 101.49 1.3125 ;
      RECT  101.905 0.8975 104.35 1.3125 ;
      RECT  104.765 0.8975 107.21 1.3125 ;
      RECT  107.625 0.8975 110.07 1.3125 ;
      RECT  110.485 0.8975 112.93 1.3125 ;
      RECT  113.345 0.8975 115.79 1.3125 ;
      RECT  116.205 0.8975 118.65 1.3125 ;
      RECT  119.065 0.8975 121.51 1.3125 ;
      RECT  121.925 0.8975 124.37 1.3125 ;
      RECT  124.785 0.8975 127.23 1.3125 ;
      RECT  127.645 0.8975 130.09 1.3125 ;
      RECT  130.505 0.8975 132.95 1.3125 ;
      RECT  133.365 0.8975 135.81 1.3125 ;
      RECT  136.225 0.8975 138.67 1.3125 ;
      RECT  139.085 0.8975 141.53 1.3125 ;
      RECT  141.945 0.8975 144.39 1.3125 ;
      RECT  144.805 0.8975 147.25 1.3125 ;
      RECT  147.665 0.8975 150.11 1.3125 ;
      RECT  150.525 0.8975 152.97 1.3125 ;
      RECT  153.385 0.8975 155.83 1.3125 ;
      RECT  156.245 0.8975 158.69 1.3125 ;
      RECT  159.105 0.8975 161.55 1.3125 ;
      RECT  64.725 1.3125 94.145 71.3625 ;
      RECT  64.725 71.3625 94.145 71.7775 ;
      RECT  64.725 71.7775 94.145 102.21 ;
      RECT  94.145 1.3125 94.56 71.3625 ;
      RECT  94.145 71.7775 94.56 102.21 ;
      RECT  94.56 1.3125 161.55 71.3625 ;
      RECT  94.56 71.7775 161.55 102.21 ;
      RECT  94.56 71.3625 94.85 71.7775 ;
      RECT  95.265 71.3625 95.555 71.7775 ;
      RECT  95.97 71.3625 96.26 71.7775 ;
      RECT  96.675 71.3625 96.965 71.7775 ;
      RECT  97.38 71.3625 97.67 71.7775 ;
      RECT  98.085 71.3625 98.375 71.7775 ;
      RECT  98.79 71.3625 99.08 71.7775 ;
      RECT  99.495 71.3625 99.785 71.7775 ;
      RECT  100.2 71.3625 100.49 71.7775 ;
      RECT  100.905 71.3625 101.195 71.7775 ;
      RECT  101.61 71.3625 101.9 71.7775 ;
      RECT  102.315 71.3625 102.605 71.7775 ;
      RECT  103.02 71.3625 103.31 71.7775 ;
      RECT  103.725 71.3625 104.015 71.7775 ;
      RECT  104.43 71.3625 104.72 71.7775 ;
      RECT  105.135 71.3625 105.425 71.7775 ;
      RECT  105.84 71.3625 106.13 71.7775 ;
      RECT  106.545 71.3625 106.835 71.7775 ;
      RECT  107.25 71.3625 107.54 71.7775 ;
      RECT  107.955 71.3625 108.245 71.7775 ;
      RECT  108.66 71.3625 108.95 71.7775 ;
      RECT  109.365 71.3625 109.655 71.7775 ;
      RECT  110.07 71.3625 110.36 71.7775 ;
      RECT  110.775 71.3625 111.065 71.7775 ;
      RECT  111.48 71.3625 111.77 71.7775 ;
      RECT  112.185 71.3625 112.475 71.7775 ;
      RECT  112.89 71.3625 113.18 71.7775 ;
      RECT  113.595 71.3625 113.885 71.7775 ;
      RECT  114.3 71.3625 114.59 71.7775 ;
      RECT  115.005 71.3625 115.295 71.7775 ;
      RECT  115.71 71.3625 116.0 71.7775 ;
      RECT  116.415 71.3625 116.705 71.7775 ;
      RECT  117.12 71.3625 117.41 71.7775 ;
      RECT  117.825 71.3625 118.115 71.7775 ;
      RECT  118.53 71.3625 118.82 71.7775 ;
      RECT  119.235 71.3625 119.525 71.7775 ;
      RECT  119.94 71.3625 120.23 71.7775 ;
      RECT  120.645 71.3625 120.935 71.7775 ;
      RECT  121.35 71.3625 121.64 71.7775 ;
      RECT  122.055 71.3625 122.345 71.7775 ;
      RECT  122.76 71.3625 123.05 71.7775 ;
      RECT  123.465 71.3625 123.755 71.7775 ;
      RECT  124.17 71.3625 124.46 71.7775 ;
      RECT  124.875 71.3625 125.165 71.7775 ;
      RECT  125.58 71.3625 125.87 71.7775 ;
      RECT  126.285 71.3625 126.575 71.7775 ;
      RECT  126.99 71.3625 127.28 71.7775 ;
      RECT  127.695 71.3625 127.985 71.7775 ;
      RECT  128.4 71.3625 128.69 71.7775 ;
      RECT  129.105 71.3625 129.395 71.7775 ;
      RECT  129.81 71.3625 130.1 71.7775 ;
      RECT  130.515 71.3625 130.805 71.7775 ;
      RECT  131.22 71.3625 131.51 71.7775 ;
      RECT  131.925 71.3625 132.215 71.7775 ;
      RECT  132.63 71.3625 132.92 71.7775 ;
      RECT  133.335 71.3625 133.625 71.7775 ;
      RECT  134.04 71.3625 134.33 71.7775 ;
      RECT  134.745 71.3625 135.035 71.7775 ;
      RECT  135.45 71.3625 135.74 71.7775 ;
      RECT  136.155 71.3625 136.445 71.7775 ;
      RECT  136.86 71.3625 137.15 71.7775 ;
      RECT  137.565 71.3625 137.855 71.7775 ;
      RECT  138.27 71.3625 138.56 71.7775 ;
      RECT  138.975 71.3625 139.265 71.7775 ;
      RECT  139.68 71.3625 139.97 71.7775 ;
      RECT  140.385 71.3625 140.675 71.7775 ;
      RECT  141.09 71.3625 141.38 71.7775 ;
      RECT  141.795 71.3625 142.085 71.7775 ;
      RECT  142.5 71.3625 142.79 71.7775 ;
      RECT  143.205 71.3625 143.495 71.7775 ;
      RECT  143.91 71.3625 144.2 71.7775 ;
      RECT  144.615 71.3625 144.905 71.7775 ;
      RECT  145.32 71.3625 145.61 71.7775 ;
      RECT  146.025 71.3625 146.315 71.7775 ;
      RECT  146.73 71.3625 147.02 71.7775 ;
      RECT  147.435 71.3625 147.725 71.7775 ;
      RECT  148.14 71.3625 148.43 71.7775 ;
      RECT  148.845 71.3625 149.135 71.7775 ;
      RECT  149.55 71.3625 149.84 71.7775 ;
      RECT  150.255 71.3625 150.545 71.7775 ;
      RECT  150.96 71.3625 151.25 71.7775 ;
      RECT  151.665 71.3625 151.955 71.7775 ;
      RECT  152.37 71.3625 152.66 71.7775 ;
      RECT  153.075 71.3625 153.365 71.7775 ;
      RECT  153.78 71.3625 154.07 71.7775 ;
      RECT  154.485 71.3625 154.775 71.7775 ;
      RECT  155.19 71.3625 155.48 71.7775 ;
      RECT  155.895 71.3625 156.185 71.7775 ;
      RECT  156.6 71.3625 156.89 71.7775 ;
      RECT  157.305 71.3625 157.595 71.7775 ;
      RECT  158.01 71.3625 158.3 71.7775 ;
      RECT  158.715 71.3625 159.005 71.7775 ;
      RECT  159.42 71.3625 159.71 71.7775 ;
      RECT  160.125 71.3625 160.415 71.7775 ;
      RECT  160.83 71.3625 161.12 71.7775 ;
      RECT  161.535 71.3625 161.55 71.7775 ;
      RECT  161.55 1.3125 161.825 71.3625 ;
      RECT  161.55 71.3625 161.825 71.7775 ;
      RECT  161.55 71.7775 161.825 127.305 ;
      RECT  161.825 1.3125 161.965 71.3625 ;
      RECT  161.825 71.7775 161.965 127.305 ;
      RECT  161.965 1.3125 162.24 71.3625 ;
      RECT  161.965 71.7775 162.24 127.305 ;
      RECT  162.24 1.3125 893.495 71.3625 ;
      RECT  162.24 71.7775 893.495 127.305 ;
      RECT  162.24 71.3625 162.53 71.7775 ;
      RECT  162.945 71.3625 163.235 71.7775 ;
      RECT  163.65 71.3625 163.94 71.7775 ;
      RECT  164.355 71.3625 164.645 71.7775 ;
      RECT  165.06 71.3625 165.35 71.7775 ;
      RECT  165.765 71.3625 166.055 71.7775 ;
      RECT  166.47 71.3625 166.76 71.7775 ;
      RECT  167.175 71.3625 167.465 71.7775 ;
      RECT  167.88 71.3625 168.17 71.7775 ;
      RECT  168.585 71.3625 168.875 71.7775 ;
      RECT  169.29 71.3625 169.58 71.7775 ;
      RECT  169.995 71.3625 170.285 71.7775 ;
      RECT  170.7 71.3625 170.99 71.7775 ;
      RECT  171.405 71.3625 171.695 71.7775 ;
      RECT  172.11 71.3625 172.4 71.7775 ;
      RECT  172.815 71.3625 173.105 71.7775 ;
      RECT  173.52 71.3625 173.81 71.7775 ;
      RECT  174.225 71.3625 174.515 71.7775 ;
      RECT  174.93 71.3625 175.22 71.7775 ;
      RECT  175.635 71.3625 175.925 71.7775 ;
      RECT  176.34 71.3625 176.63 71.7775 ;
      RECT  177.045 71.3625 177.335 71.7775 ;
      RECT  177.75 71.3625 178.04 71.7775 ;
      RECT  178.455 71.3625 178.745 71.7775 ;
      RECT  179.16 71.3625 179.45 71.7775 ;
      RECT  179.865 71.3625 180.155 71.7775 ;
      RECT  180.57 71.3625 180.86 71.7775 ;
      RECT  181.275 71.3625 181.565 71.7775 ;
      RECT  181.98 71.3625 182.27 71.7775 ;
      RECT  182.685 71.3625 182.975 71.7775 ;
      RECT  183.39 71.3625 183.68 71.7775 ;
      RECT  184.095 71.3625 184.385 71.7775 ;
      RECT  184.8 71.3625 185.09 71.7775 ;
      RECT  185.505 71.3625 185.795 71.7775 ;
      RECT  186.21 71.3625 186.5 71.7775 ;
      RECT  186.915 71.3625 187.205 71.7775 ;
      RECT  187.62 71.3625 187.91 71.7775 ;
      RECT  188.325 71.3625 188.615 71.7775 ;
      RECT  189.03 71.3625 189.32 71.7775 ;
      RECT  189.735 71.3625 190.025 71.7775 ;
      RECT  190.44 71.3625 190.73 71.7775 ;
      RECT  191.145 71.3625 191.435 71.7775 ;
      RECT  191.85 71.3625 192.14 71.7775 ;
      RECT  192.555 71.3625 192.845 71.7775 ;
      RECT  193.26 71.3625 193.55 71.7775 ;
      RECT  193.965 71.3625 194.255 71.7775 ;
      RECT  194.67 71.3625 194.96 71.7775 ;
      RECT  195.375 71.3625 195.665 71.7775 ;
      RECT  196.08 71.3625 196.37 71.7775 ;
      RECT  196.785 71.3625 197.075 71.7775 ;
      RECT  197.49 71.3625 197.78 71.7775 ;
      RECT  198.195 71.3625 198.485 71.7775 ;
      RECT  198.9 71.3625 199.19 71.7775 ;
      RECT  199.605 71.3625 199.895 71.7775 ;
      RECT  200.31 71.3625 200.6 71.7775 ;
      RECT  201.015 71.3625 201.305 71.7775 ;
      RECT  201.72 71.3625 202.01 71.7775 ;
      RECT  202.425 71.3625 202.715 71.7775 ;
      RECT  203.13 71.3625 203.42 71.7775 ;
      RECT  203.835 71.3625 204.125 71.7775 ;
      RECT  204.54 71.3625 204.83 71.7775 ;
      RECT  205.245 71.3625 205.535 71.7775 ;
      RECT  205.95 71.3625 206.24 71.7775 ;
      RECT  206.655 71.3625 206.945 71.7775 ;
      RECT  207.36 71.3625 207.65 71.7775 ;
      RECT  208.065 71.3625 208.355 71.7775 ;
      RECT  208.77 71.3625 209.06 71.7775 ;
      RECT  209.475 71.3625 209.765 71.7775 ;
      RECT  210.18 71.3625 210.47 71.7775 ;
      RECT  210.885 71.3625 211.175 71.7775 ;
      RECT  211.59 71.3625 211.88 71.7775 ;
      RECT  212.295 71.3625 212.585 71.7775 ;
      RECT  213.0 71.3625 213.29 71.7775 ;
      RECT  213.705 71.3625 213.995 71.7775 ;
      RECT  214.41 71.3625 214.7 71.7775 ;
      RECT  215.115 71.3625 215.405 71.7775 ;
      RECT  215.82 71.3625 216.11 71.7775 ;
      RECT  216.525 71.3625 216.815 71.7775 ;
      RECT  217.23 71.3625 217.52 71.7775 ;
      RECT  217.935 71.3625 218.225 71.7775 ;
      RECT  218.64 71.3625 218.93 71.7775 ;
      RECT  219.345 71.3625 219.635 71.7775 ;
      RECT  220.05 71.3625 220.34 71.7775 ;
      RECT  220.755 71.3625 221.045 71.7775 ;
      RECT  221.46 71.3625 221.75 71.7775 ;
      RECT  222.165 71.3625 222.455 71.7775 ;
      RECT  222.87 71.3625 223.16 71.7775 ;
      RECT  223.575 71.3625 223.865 71.7775 ;
      RECT  224.28 71.3625 224.57 71.7775 ;
      RECT  224.985 71.3625 225.275 71.7775 ;
      RECT  225.69 71.3625 225.98 71.7775 ;
      RECT  226.395 71.3625 226.685 71.7775 ;
      RECT  227.1 71.3625 227.39 71.7775 ;
      RECT  227.805 71.3625 228.095 71.7775 ;
      RECT  228.51 71.3625 228.8 71.7775 ;
      RECT  229.215 71.3625 229.505 71.7775 ;
      RECT  229.92 71.3625 230.21 71.7775 ;
      RECT  230.625 71.3625 230.915 71.7775 ;
      RECT  231.33 71.3625 231.62 71.7775 ;
      RECT  232.035 71.3625 232.325 71.7775 ;
      RECT  232.74 71.3625 233.03 71.7775 ;
      RECT  233.445 71.3625 233.735 71.7775 ;
      RECT  234.15 71.3625 234.44 71.7775 ;
      RECT  234.855 71.3625 235.145 71.7775 ;
      RECT  235.56 71.3625 235.85 71.7775 ;
      RECT  236.265 71.3625 236.555 71.7775 ;
      RECT  236.97 71.3625 237.26 71.7775 ;
      RECT  237.675 71.3625 237.965 71.7775 ;
      RECT  238.38 71.3625 238.67 71.7775 ;
      RECT  239.085 71.3625 239.375 71.7775 ;
      RECT  239.79 71.3625 240.08 71.7775 ;
      RECT  240.495 71.3625 240.785 71.7775 ;
      RECT  241.2 71.3625 241.49 71.7775 ;
      RECT  241.905 71.3625 242.195 71.7775 ;
      RECT  242.61 71.3625 242.9 71.7775 ;
      RECT  243.315 71.3625 243.605 71.7775 ;
      RECT  244.02 71.3625 244.31 71.7775 ;
      RECT  244.725 71.3625 245.015 71.7775 ;
      RECT  245.43 71.3625 245.72 71.7775 ;
      RECT  246.135 71.3625 246.425 71.7775 ;
      RECT  246.84 71.3625 247.13 71.7775 ;
      RECT  247.545 71.3625 247.835 71.7775 ;
      RECT  248.25 71.3625 248.54 71.7775 ;
      RECT  248.955 71.3625 249.245 71.7775 ;
      RECT  249.66 71.3625 249.95 71.7775 ;
      RECT  250.365 71.3625 250.655 71.7775 ;
      RECT  251.07 71.3625 251.36 71.7775 ;
      RECT  251.775 71.3625 252.065 71.7775 ;
      RECT  252.48 71.3625 252.77 71.7775 ;
      RECT  253.185 71.3625 253.475 71.7775 ;
      RECT  253.89 71.3625 254.18 71.7775 ;
      RECT  254.595 71.3625 254.885 71.7775 ;
      RECT  255.3 71.3625 255.59 71.7775 ;
      RECT  256.005 71.3625 256.295 71.7775 ;
      RECT  256.71 71.3625 257.0 71.7775 ;
      RECT  257.415 71.3625 257.705 71.7775 ;
      RECT  258.12 71.3625 258.41 71.7775 ;
      RECT  258.825 71.3625 259.115 71.7775 ;
      RECT  259.53 71.3625 259.82 71.7775 ;
      RECT  260.235 71.3625 260.525 71.7775 ;
      RECT  260.94 71.3625 261.23 71.7775 ;
      RECT  261.645 71.3625 261.935 71.7775 ;
      RECT  262.35 71.3625 262.64 71.7775 ;
      RECT  263.055 71.3625 263.345 71.7775 ;
      RECT  263.76 71.3625 264.05 71.7775 ;
      RECT  264.465 71.3625 264.755 71.7775 ;
      RECT  265.17 71.3625 265.46 71.7775 ;
      RECT  265.875 71.3625 266.165 71.7775 ;
      RECT  266.58 71.3625 266.87 71.7775 ;
      RECT  267.285 71.3625 267.575 71.7775 ;
      RECT  267.99 71.3625 268.28 71.7775 ;
      RECT  268.695 71.3625 268.985 71.7775 ;
      RECT  269.4 71.3625 269.69 71.7775 ;
      RECT  270.105 71.3625 270.395 71.7775 ;
      RECT  270.81 71.3625 271.1 71.7775 ;
      RECT  271.515 71.3625 271.805 71.7775 ;
      RECT  272.22 71.3625 272.51 71.7775 ;
      RECT  272.925 71.3625 273.215 71.7775 ;
      RECT  273.63 71.3625 273.92 71.7775 ;
      RECT  274.335 71.3625 893.495 71.7775 ;
   LAYER  metal4 ;
      RECT  0.14 0.14 893.495 127.305 ;
   END
END    mp3_data_array_2
END    LIBRARY
