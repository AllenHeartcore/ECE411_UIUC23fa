VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO mp3_tag_array_2
   CLASS BLOCK ;
   SIZE 84.86 BY 48.055 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  22.155 1.0375 22.29 1.1725 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  25.015 1.0375 25.15 1.1725 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  27.875 1.0375 28.01 1.1725 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  30.735 1.0375 30.87 1.1725 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  33.595 1.0375 33.73 1.1725 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.455 1.0375 36.59 1.1725 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  39.315 1.0375 39.45 1.1725 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  42.175 1.0375 42.31 1.1725 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.035 1.0375 45.17 1.1725 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.895 1.0375 48.03 1.1725 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  50.755 1.0375 50.89 1.1725 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  53.615 1.0375 53.75 1.1725 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.475 1.0375 56.61 1.1725 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.335 1.0375 59.47 1.1725 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  62.195 1.0375 62.33 1.1725 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  65.055 1.0375 65.19 1.1725 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.915 1.0375 68.05 1.1725 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.775 1.0375 70.91 1.1725 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.635 1.0375 73.77 1.1725 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.495 1.0375 76.63 1.1725 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  79.355 1.0375 79.49 1.1725 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.215 1.0375 82.35 1.1725 ;
      END
   END din0[21]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  19.295 1.0375 19.43 1.1725 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.575 39.2125 13.71 39.3475 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.575 41.9425 13.71 42.0775 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.575 44.1525 13.71 44.2875 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.575 46.8825 13.71 47.0175 ;
      END
   END addr0[4]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 2.6825 0.42 2.8175 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 5.4125 0.42 5.5475 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.5275 2.7675 6.6625 2.9025 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  31.495 10.87 31.63 11.005 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.905 10.87 33.04 11.005 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  34.315 10.87 34.45 11.005 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.725 10.87 35.86 11.005 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.135 10.87 37.27 11.005 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  38.545 10.87 38.68 11.005 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  39.955 10.87 40.09 11.005 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  41.365 10.87 41.5 11.005 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  42.775 10.87 42.91 11.005 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  44.185 10.87 44.32 11.005 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.595 10.87 45.73 11.005 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.005 10.87 47.14 11.005 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  48.415 10.87 48.55 11.005 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  49.825 10.87 49.96 11.005 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  51.235 10.87 51.37 11.005 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.645 10.87 52.78 11.005 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  54.055 10.87 54.19 11.005 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.465 10.87 55.6 11.005 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.875 10.87 57.01 11.005 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  58.285 10.87 58.42 11.005 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.695 10.87 59.83 11.005 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.105 10.87 61.24 11.005 ;
      END
   END dout0[21]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 84.72 47.915 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 84.72 47.915 ;
   LAYER  metal3 ;
      RECT  0.14 0.14 22.015 0.8975 ;
      RECT  22.015 0.14 22.43 0.8975 ;
      RECT  22.015 1.3125 22.43 47.915 ;
      RECT  22.43 0.14 84.72 0.8975 ;
      RECT  22.43 0.8975 24.875 1.3125 ;
      RECT  25.29 0.8975 27.735 1.3125 ;
      RECT  28.15 0.8975 30.595 1.3125 ;
      RECT  31.01 0.8975 33.455 1.3125 ;
      RECT  33.87 0.8975 36.315 1.3125 ;
      RECT  36.73 0.8975 39.175 1.3125 ;
      RECT  39.59 0.8975 42.035 1.3125 ;
      RECT  42.45 0.8975 44.895 1.3125 ;
      RECT  45.31 0.8975 47.755 1.3125 ;
      RECT  48.17 0.8975 50.615 1.3125 ;
      RECT  51.03 0.8975 53.475 1.3125 ;
      RECT  53.89 0.8975 56.335 1.3125 ;
      RECT  56.75 0.8975 59.195 1.3125 ;
      RECT  59.61 0.8975 62.055 1.3125 ;
      RECT  62.47 0.8975 64.915 1.3125 ;
      RECT  65.33 0.8975 67.775 1.3125 ;
      RECT  68.19 0.8975 70.635 1.3125 ;
      RECT  71.05 0.8975 73.495 1.3125 ;
      RECT  73.91 0.8975 76.355 1.3125 ;
      RECT  76.77 0.8975 79.215 1.3125 ;
      RECT  79.63 0.8975 82.075 1.3125 ;
      RECT  82.49 0.8975 84.72 1.3125 ;
      RECT  0.14 0.8975 19.155 1.3125 ;
      RECT  19.57 0.8975 22.015 1.3125 ;
      RECT  0.14 39.0725 13.435 39.4875 ;
      RECT  0.14 39.4875 13.435 47.915 ;
      RECT  13.435 1.3125 13.85 39.0725 ;
      RECT  13.85 1.3125 22.015 39.0725 ;
      RECT  13.85 39.0725 22.015 39.4875 ;
      RECT  13.85 39.4875 22.015 47.915 ;
      RECT  13.435 39.4875 13.85 41.8025 ;
      RECT  13.435 42.2175 13.85 44.0125 ;
      RECT  13.435 44.4275 13.85 46.7425 ;
      RECT  13.435 47.1575 13.85 47.915 ;
      RECT  0.14 1.3125 0.145 2.5425 ;
      RECT  0.14 2.5425 0.145 2.9575 ;
      RECT  0.14 2.9575 0.145 39.0725 ;
      RECT  0.145 1.3125 0.56 2.5425 ;
      RECT  0.56 1.3125 13.435 2.5425 ;
      RECT  0.145 2.9575 0.56 5.2725 ;
      RECT  0.145 5.6875 0.56 39.0725 ;
      RECT  0.56 2.5425 6.3875 2.6275 ;
      RECT  0.56 2.6275 6.3875 2.9575 ;
      RECT  6.3875 2.5425 6.8025 2.6275 ;
      RECT  6.8025 2.5425 13.435 2.6275 ;
      RECT  6.8025 2.6275 13.435 2.9575 ;
      RECT  0.56 2.9575 6.3875 3.0425 ;
      RECT  0.56 3.0425 6.3875 39.0725 ;
      RECT  6.3875 3.0425 6.8025 39.0725 ;
      RECT  6.8025 2.9575 13.435 3.0425 ;
      RECT  6.8025 3.0425 13.435 39.0725 ;
      RECT  22.43 1.3125 31.355 10.73 ;
      RECT  22.43 10.73 31.355 11.145 ;
      RECT  22.43 11.145 31.355 47.915 ;
      RECT  31.355 1.3125 31.77 10.73 ;
      RECT  31.355 11.145 31.77 47.915 ;
      RECT  31.77 1.3125 84.72 10.73 ;
      RECT  31.77 11.145 84.72 47.915 ;
      RECT  31.77 10.73 32.765 11.145 ;
      RECT  33.18 10.73 34.175 11.145 ;
      RECT  34.59 10.73 35.585 11.145 ;
      RECT  36.0 10.73 36.995 11.145 ;
      RECT  37.41 10.73 38.405 11.145 ;
      RECT  38.82 10.73 39.815 11.145 ;
      RECT  40.23 10.73 41.225 11.145 ;
      RECT  41.64 10.73 42.635 11.145 ;
      RECT  43.05 10.73 44.045 11.145 ;
      RECT  44.46 10.73 45.455 11.145 ;
      RECT  45.87 10.73 46.865 11.145 ;
      RECT  47.28 10.73 48.275 11.145 ;
      RECT  48.69 10.73 49.685 11.145 ;
      RECT  50.1 10.73 51.095 11.145 ;
      RECT  51.51 10.73 52.505 11.145 ;
      RECT  52.92 10.73 53.915 11.145 ;
      RECT  54.33 10.73 55.325 11.145 ;
      RECT  55.74 10.73 56.735 11.145 ;
      RECT  57.15 10.73 58.145 11.145 ;
      RECT  58.56 10.73 59.555 11.145 ;
      RECT  59.97 10.73 60.965 11.145 ;
      RECT  61.38 10.73 84.72 11.145 ;
   LAYER  metal4 ;
      RECT  0.14 0.14 84.72 47.915 ;
   END
END    mp3_tag_array_2
END    LIBRARY
