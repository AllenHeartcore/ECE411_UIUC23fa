VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO mp3_tag_array_1
   CLASS BLOCK ;
   SIZE 87.72 BY 46.78 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  19.295 1.0375 19.43 1.1725 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  22.155 1.0375 22.29 1.1725 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  25.015 1.0375 25.15 1.1725 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  27.875 1.0375 28.01 1.1725 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  30.735 1.0375 30.87 1.1725 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  33.595 1.0375 33.73 1.1725 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.455 1.0375 36.59 1.1725 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  39.315 1.0375 39.45 1.1725 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  42.175 1.0375 42.31 1.1725 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.035 1.0375 45.17 1.1725 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.895 1.0375 48.03 1.1725 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  50.755 1.0375 50.89 1.1725 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  53.615 1.0375 53.75 1.1725 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.475 1.0375 56.61 1.1725 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.335 1.0375 59.47 1.1725 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  62.195 1.0375 62.33 1.1725 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  65.055 1.0375 65.19 1.1725 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.915 1.0375 68.05 1.1725 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.775 1.0375 70.91 1.1725 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.635 1.0375 73.77 1.1725 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.495 1.0375 76.63 1.1725 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  79.355 1.0375 79.49 1.1725 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.215 1.0375 82.35 1.1725 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.075 1.0375 85.21 1.1725 ;
      END
   END din0[23]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.575 37.9375 13.71 38.0725 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.575 40.6675 13.71 40.8025 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.575 42.8775 13.71 43.0125 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.575 45.6075 13.71 45.7425 ;
      END
   END addr0[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 1.4075 0.42 1.5425 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 4.1375 0.42 4.2725 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.5275 1.4925 6.6625 1.6275 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  30.395 12.55 30.53 12.685 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  31.1 12.55 31.235 12.685 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  31.805 12.55 31.94 12.685 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.51 12.55 32.645 12.685 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  33.215 12.55 33.35 12.685 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  33.92 12.55 34.055 12.685 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  34.625 12.55 34.76 12.685 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.33 12.55 35.465 12.685 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.035 12.55 36.17 12.685 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.74 12.55 36.875 12.685 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.445 12.55 37.58 12.685 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  38.15 12.55 38.285 12.685 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  38.855 12.55 38.99 12.685 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  39.56 12.55 39.695 12.685 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.265 12.55 40.4 12.685 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.97 12.55 41.105 12.685 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  41.675 12.55 41.81 12.685 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  42.38 12.55 42.515 12.685 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.085 12.55 43.22 12.685 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.79 12.55 43.925 12.685 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  44.495 12.55 44.63 12.685 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.2 12.55 45.335 12.685 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.905 12.55 46.04 12.685 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  46.61 12.55 46.745 12.685 ;
      END
   END dout0[23]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 87.58 46.64 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 87.58 46.64 ;
   LAYER  metal3 ;
      RECT  0.14 0.14 19.155 0.8975 ;
      RECT  19.155 0.14 19.57 0.8975 ;
      RECT  19.155 1.3125 19.57 46.64 ;
      RECT  19.57 0.14 87.58 0.8975 ;
      RECT  19.57 0.8975 22.015 1.3125 ;
      RECT  22.43 0.8975 24.875 1.3125 ;
      RECT  25.29 0.8975 27.735 1.3125 ;
      RECT  28.15 0.8975 30.595 1.3125 ;
      RECT  31.01 0.8975 33.455 1.3125 ;
      RECT  33.87 0.8975 36.315 1.3125 ;
      RECT  36.73 0.8975 39.175 1.3125 ;
      RECT  39.59 0.8975 42.035 1.3125 ;
      RECT  42.45 0.8975 44.895 1.3125 ;
      RECT  45.31 0.8975 47.755 1.3125 ;
      RECT  48.17 0.8975 50.615 1.3125 ;
      RECT  51.03 0.8975 53.475 1.3125 ;
      RECT  53.89 0.8975 56.335 1.3125 ;
      RECT  56.75 0.8975 59.195 1.3125 ;
      RECT  59.61 0.8975 62.055 1.3125 ;
      RECT  62.47 0.8975 64.915 1.3125 ;
      RECT  65.33 0.8975 67.775 1.3125 ;
      RECT  68.19 0.8975 70.635 1.3125 ;
      RECT  71.05 0.8975 73.495 1.3125 ;
      RECT  73.91 0.8975 76.355 1.3125 ;
      RECT  76.77 0.8975 79.215 1.3125 ;
      RECT  79.63 0.8975 82.075 1.3125 ;
      RECT  82.49 0.8975 84.935 1.3125 ;
      RECT  85.35 0.8975 87.58 1.3125 ;
      RECT  0.14 37.7975 13.435 38.2125 ;
      RECT  0.14 38.2125 13.435 46.64 ;
      RECT  13.435 1.3125 13.85 37.7975 ;
      RECT  13.85 1.3125 19.155 37.7975 ;
      RECT  13.85 37.7975 19.155 38.2125 ;
      RECT  13.85 38.2125 19.155 46.64 ;
      RECT  13.435 38.2125 13.85 40.5275 ;
      RECT  13.435 40.9425 13.85 42.7375 ;
      RECT  13.435 43.1525 13.85 45.4675 ;
      RECT  13.435 45.8825 13.85 46.64 ;
      RECT  0.14 0.8975 0.145 1.2675 ;
      RECT  0.14 1.2675 0.145 1.3125 ;
      RECT  0.145 0.8975 0.56 1.2675 ;
      RECT  0.56 0.8975 19.155 1.2675 ;
      RECT  0.56 1.2675 19.155 1.3125 ;
      RECT  0.14 1.3125 0.145 1.6825 ;
      RECT  0.14 1.6825 0.145 37.7975 ;
      RECT  0.145 1.6825 0.56 3.9975 ;
      RECT  0.145 4.4125 0.56 37.7975 ;
      RECT  0.56 1.3125 6.3875 1.3525 ;
      RECT  0.56 1.3525 6.3875 1.6825 ;
      RECT  6.3875 1.3125 6.8025 1.3525 ;
      RECT  6.8025 1.3125 13.435 1.3525 ;
      RECT  6.8025 1.3525 13.435 1.6825 ;
      RECT  0.56 1.6825 6.3875 1.7675 ;
      RECT  0.56 1.7675 6.3875 37.7975 ;
      RECT  6.3875 1.7675 6.8025 37.7975 ;
      RECT  6.8025 1.6825 13.435 1.7675 ;
      RECT  6.8025 1.7675 13.435 37.7975 ;
      RECT  19.57 1.3125 30.255 12.41 ;
      RECT  19.57 12.41 30.255 12.825 ;
      RECT  19.57 12.825 30.255 46.64 ;
      RECT  30.255 1.3125 30.67 12.41 ;
      RECT  30.255 12.825 30.67 46.64 ;
      RECT  30.67 1.3125 87.58 12.41 ;
      RECT  30.67 12.825 87.58 46.64 ;
      RECT  30.67 12.41 30.96 12.825 ;
      RECT  31.375 12.41 31.665 12.825 ;
      RECT  32.08 12.41 32.37 12.825 ;
      RECT  32.785 12.41 33.075 12.825 ;
      RECT  33.49 12.41 33.78 12.825 ;
      RECT  34.195 12.41 34.485 12.825 ;
      RECT  34.9 12.41 35.19 12.825 ;
      RECT  35.605 12.41 35.895 12.825 ;
      RECT  36.31 12.41 36.6 12.825 ;
      RECT  37.015 12.41 37.305 12.825 ;
      RECT  37.72 12.41 38.01 12.825 ;
      RECT  38.425 12.41 38.715 12.825 ;
      RECT  39.13 12.41 39.42 12.825 ;
      RECT  39.835 12.41 40.125 12.825 ;
      RECT  40.54 12.41 40.83 12.825 ;
      RECT  41.245 12.41 41.535 12.825 ;
      RECT  41.95 12.41 42.24 12.825 ;
      RECT  42.655 12.41 42.945 12.825 ;
      RECT  43.36 12.41 43.65 12.825 ;
      RECT  44.065 12.41 44.355 12.825 ;
      RECT  44.77 12.41 45.06 12.825 ;
      RECT  45.475 12.41 45.765 12.825 ;
      RECT  46.18 12.41 46.47 12.825 ;
      RECT  46.885 12.41 87.58 12.825 ;
   LAYER  metal4 ;
      RECT  0.14 0.14 87.58 46.64 ;
   END
END    mp3_tag_array_1
END    LIBRARY
