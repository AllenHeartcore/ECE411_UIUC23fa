VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO mp3_data_array
   CLASS BLOCK ;
   SIZE 893.36 BY 125.11 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  161.415 1.0375 161.55 1.1725 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  164.275 1.0375 164.41 1.1725 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  167.135 1.0375 167.27 1.1725 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.995 1.0375 170.13 1.1725 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.855 1.0375 172.99 1.1725 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  175.715 1.0375 175.85 1.1725 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.575 1.0375 178.71 1.1725 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  181.435 1.0375 181.57 1.1725 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  184.295 1.0375 184.43 1.1725 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  187.155 1.0375 187.29 1.1725 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  190.015 1.0375 190.15 1.1725 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.875 1.0375 193.01 1.1725 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  195.735 1.0375 195.87 1.1725 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  198.595 1.0375 198.73 1.1725 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  201.455 1.0375 201.59 1.1725 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  204.315 1.0375 204.45 1.1725 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  207.175 1.0375 207.31 1.1725 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  210.035 1.0375 210.17 1.1725 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.895 1.0375 213.03 1.1725 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  215.755 1.0375 215.89 1.1725 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  218.615 1.0375 218.75 1.1725 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  221.475 1.0375 221.61 1.1725 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  224.335 1.0375 224.47 1.1725 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  227.195 1.0375 227.33 1.1725 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  230.055 1.0375 230.19 1.1725 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  232.915 1.0375 233.05 1.1725 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  235.775 1.0375 235.91 1.1725 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  238.635 1.0375 238.77 1.1725 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  241.495 1.0375 241.63 1.1725 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  244.355 1.0375 244.49 1.1725 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  247.215 1.0375 247.35 1.1725 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  250.075 1.0375 250.21 1.1725 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  252.935 1.0375 253.07 1.1725 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  255.795 1.0375 255.93 1.1725 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  258.655 1.0375 258.79 1.1725 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  261.515 1.0375 261.65 1.1725 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  264.375 1.0375 264.51 1.1725 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  267.235 1.0375 267.37 1.1725 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  270.095 1.0375 270.23 1.1725 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  272.955 1.0375 273.09 1.1725 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  275.815 1.0375 275.95 1.1725 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  278.675 1.0375 278.81 1.1725 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  281.535 1.0375 281.67 1.1725 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  284.395 1.0375 284.53 1.1725 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  287.255 1.0375 287.39 1.1725 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  290.115 1.0375 290.25 1.1725 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  292.975 1.0375 293.11 1.1725 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  295.835 1.0375 295.97 1.1725 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  298.695 1.0375 298.83 1.1725 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  301.555 1.0375 301.69 1.1725 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  304.415 1.0375 304.55 1.1725 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  307.275 1.0375 307.41 1.1725 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  310.135 1.0375 310.27 1.1725 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  312.995 1.0375 313.13 1.1725 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  315.855 1.0375 315.99 1.1725 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  318.715 1.0375 318.85 1.1725 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  321.575 1.0375 321.71 1.1725 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  324.435 1.0375 324.57 1.1725 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  327.295 1.0375 327.43 1.1725 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  330.155 1.0375 330.29 1.1725 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  333.015 1.0375 333.15 1.1725 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  335.875 1.0375 336.01 1.1725 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  338.735 1.0375 338.87 1.1725 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  341.595 1.0375 341.73 1.1725 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  344.455 1.0375 344.59 1.1725 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  347.315 1.0375 347.45 1.1725 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  350.175 1.0375 350.31 1.1725 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  353.035 1.0375 353.17 1.1725 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  355.895 1.0375 356.03 1.1725 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  358.755 1.0375 358.89 1.1725 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  361.615 1.0375 361.75 1.1725 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  364.475 1.0375 364.61 1.1725 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  367.335 1.0375 367.47 1.1725 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  370.195 1.0375 370.33 1.1725 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  373.055 1.0375 373.19 1.1725 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  375.915 1.0375 376.05 1.1725 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  378.775 1.0375 378.91 1.1725 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  381.635 1.0375 381.77 1.1725 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  384.495 1.0375 384.63 1.1725 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  387.355 1.0375 387.49 1.1725 ;
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  390.215 1.0375 390.35 1.1725 ;
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  393.075 1.0375 393.21 1.1725 ;
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  395.935 1.0375 396.07 1.1725 ;
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  398.795 1.0375 398.93 1.1725 ;
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  401.655 1.0375 401.79 1.1725 ;
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  404.515 1.0375 404.65 1.1725 ;
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  407.375 1.0375 407.51 1.1725 ;
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  410.235 1.0375 410.37 1.1725 ;
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  413.095 1.0375 413.23 1.1725 ;
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  415.955 1.0375 416.09 1.1725 ;
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  418.815 1.0375 418.95 1.1725 ;
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  421.675 1.0375 421.81 1.1725 ;
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  424.535 1.0375 424.67 1.1725 ;
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  427.395 1.0375 427.53 1.1725 ;
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  430.255 1.0375 430.39 1.1725 ;
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  433.115 1.0375 433.25 1.1725 ;
      END
   END din0[95]
   PIN din0[96]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  435.975 1.0375 436.11 1.1725 ;
      END
   END din0[96]
   PIN din0[97]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  438.835 1.0375 438.97 1.1725 ;
      END
   END din0[97]
   PIN din0[98]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  441.695 1.0375 441.83 1.1725 ;
      END
   END din0[98]
   PIN din0[99]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  444.555 1.0375 444.69 1.1725 ;
      END
   END din0[99]
   PIN din0[100]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  447.415 1.0375 447.55 1.1725 ;
      END
   END din0[100]
   PIN din0[101]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  450.275 1.0375 450.41 1.1725 ;
      END
   END din0[101]
   PIN din0[102]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  453.135 1.0375 453.27 1.1725 ;
      END
   END din0[102]
   PIN din0[103]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  455.995 1.0375 456.13 1.1725 ;
      END
   END din0[103]
   PIN din0[104]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  458.855 1.0375 458.99 1.1725 ;
      END
   END din0[104]
   PIN din0[105]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  461.715 1.0375 461.85 1.1725 ;
      END
   END din0[105]
   PIN din0[106]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  464.575 1.0375 464.71 1.1725 ;
      END
   END din0[106]
   PIN din0[107]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  467.435 1.0375 467.57 1.1725 ;
      END
   END din0[107]
   PIN din0[108]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  470.295 1.0375 470.43 1.1725 ;
      END
   END din0[108]
   PIN din0[109]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  473.155 1.0375 473.29 1.1725 ;
      END
   END din0[109]
   PIN din0[110]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  476.015 1.0375 476.15 1.1725 ;
      END
   END din0[110]
   PIN din0[111]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  478.875 1.0375 479.01 1.1725 ;
      END
   END din0[111]
   PIN din0[112]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  481.735 1.0375 481.87 1.1725 ;
      END
   END din0[112]
   PIN din0[113]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  484.595 1.0375 484.73 1.1725 ;
      END
   END din0[113]
   PIN din0[114]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  487.455 1.0375 487.59 1.1725 ;
      END
   END din0[114]
   PIN din0[115]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  490.315 1.0375 490.45 1.1725 ;
      END
   END din0[115]
   PIN din0[116]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  493.175 1.0375 493.31 1.1725 ;
      END
   END din0[116]
   PIN din0[117]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  496.035 1.0375 496.17 1.1725 ;
      END
   END din0[117]
   PIN din0[118]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  498.895 1.0375 499.03 1.1725 ;
      END
   END din0[118]
   PIN din0[119]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  501.755 1.0375 501.89 1.1725 ;
      END
   END din0[119]
   PIN din0[120]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  504.615 1.0375 504.75 1.1725 ;
      END
   END din0[120]
   PIN din0[121]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  507.475 1.0375 507.61 1.1725 ;
      END
   END din0[121]
   PIN din0[122]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  510.335 1.0375 510.47 1.1725 ;
      END
   END din0[122]
   PIN din0[123]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  513.195 1.0375 513.33 1.1725 ;
      END
   END din0[123]
   PIN din0[124]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  516.055 1.0375 516.19 1.1725 ;
      END
   END din0[124]
   PIN din0[125]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  518.915 1.0375 519.05 1.1725 ;
      END
   END din0[125]
   PIN din0[126]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  521.775 1.0375 521.91 1.1725 ;
      END
   END din0[126]
   PIN din0[127]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  524.635 1.0375 524.77 1.1725 ;
      END
   END din0[127]
   PIN din0[128]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  527.495 1.0375 527.63 1.1725 ;
      END
   END din0[128]
   PIN din0[129]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  530.355 1.0375 530.49 1.1725 ;
      END
   END din0[129]
   PIN din0[130]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  533.215 1.0375 533.35 1.1725 ;
      END
   END din0[130]
   PIN din0[131]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  536.075 1.0375 536.21 1.1725 ;
      END
   END din0[131]
   PIN din0[132]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  538.935 1.0375 539.07 1.1725 ;
      END
   END din0[132]
   PIN din0[133]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  541.795 1.0375 541.93 1.1725 ;
      END
   END din0[133]
   PIN din0[134]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  544.655 1.0375 544.79 1.1725 ;
      END
   END din0[134]
   PIN din0[135]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  547.515 1.0375 547.65 1.1725 ;
      END
   END din0[135]
   PIN din0[136]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  550.375 1.0375 550.51 1.1725 ;
      END
   END din0[136]
   PIN din0[137]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  553.235 1.0375 553.37 1.1725 ;
      END
   END din0[137]
   PIN din0[138]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  556.095 1.0375 556.23 1.1725 ;
      END
   END din0[138]
   PIN din0[139]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  558.955 1.0375 559.09 1.1725 ;
      END
   END din0[139]
   PIN din0[140]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  561.815 1.0375 561.95 1.1725 ;
      END
   END din0[140]
   PIN din0[141]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  564.675 1.0375 564.81 1.1725 ;
      END
   END din0[141]
   PIN din0[142]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  567.535 1.0375 567.67 1.1725 ;
      END
   END din0[142]
   PIN din0[143]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  570.395 1.0375 570.53 1.1725 ;
      END
   END din0[143]
   PIN din0[144]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  573.255 1.0375 573.39 1.1725 ;
      END
   END din0[144]
   PIN din0[145]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  576.115 1.0375 576.25 1.1725 ;
      END
   END din0[145]
   PIN din0[146]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  578.975 1.0375 579.11 1.1725 ;
      END
   END din0[146]
   PIN din0[147]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  581.835 1.0375 581.97 1.1725 ;
      END
   END din0[147]
   PIN din0[148]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  584.695 1.0375 584.83 1.1725 ;
      END
   END din0[148]
   PIN din0[149]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  587.555 1.0375 587.69 1.1725 ;
      END
   END din0[149]
   PIN din0[150]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  590.415 1.0375 590.55 1.1725 ;
      END
   END din0[150]
   PIN din0[151]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  593.275 1.0375 593.41 1.1725 ;
      END
   END din0[151]
   PIN din0[152]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  596.135 1.0375 596.27 1.1725 ;
      END
   END din0[152]
   PIN din0[153]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  598.995 1.0375 599.13 1.1725 ;
      END
   END din0[153]
   PIN din0[154]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  601.855 1.0375 601.99 1.1725 ;
      END
   END din0[154]
   PIN din0[155]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  604.715 1.0375 604.85 1.1725 ;
      END
   END din0[155]
   PIN din0[156]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  607.575 1.0375 607.71 1.1725 ;
      END
   END din0[156]
   PIN din0[157]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  610.435 1.0375 610.57 1.1725 ;
      END
   END din0[157]
   PIN din0[158]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  613.295 1.0375 613.43 1.1725 ;
      END
   END din0[158]
   PIN din0[159]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  616.155 1.0375 616.29 1.1725 ;
      END
   END din0[159]
   PIN din0[160]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  619.015 1.0375 619.15 1.1725 ;
      END
   END din0[160]
   PIN din0[161]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  621.875 1.0375 622.01 1.1725 ;
      END
   END din0[161]
   PIN din0[162]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  624.735 1.0375 624.87 1.1725 ;
      END
   END din0[162]
   PIN din0[163]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  627.595 1.0375 627.73 1.1725 ;
      END
   END din0[163]
   PIN din0[164]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  630.455 1.0375 630.59 1.1725 ;
      END
   END din0[164]
   PIN din0[165]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  633.315 1.0375 633.45 1.1725 ;
      END
   END din0[165]
   PIN din0[166]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  636.175 1.0375 636.31 1.1725 ;
      END
   END din0[166]
   PIN din0[167]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  639.035 1.0375 639.17 1.1725 ;
      END
   END din0[167]
   PIN din0[168]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  641.895 1.0375 642.03 1.1725 ;
      END
   END din0[168]
   PIN din0[169]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  644.755 1.0375 644.89 1.1725 ;
      END
   END din0[169]
   PIN din0[170]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  647.615 1.0375 647.75 1.1725 ;
      END
   END din0[170]
   PIN din0[171]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  650.475 1.0375 650.61 1.1725 ;
      END
   END din0[171]
   PIN din0[172]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  653.335 1.0375 653.47 1.1725 ;
      END
   END din0[172]
   PIN din0[173]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  656.195 1.0375 656.33 1.1725 ;
      END
   END din0[173]
   PIN din0[174]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  659.055 1.0375 659.19 1.1725 ;
      END
   END din0[174]
   PIN din0[175]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  661.915 1.0375 662.05 1.1725 ;
      END
   END din0[175]
   PIN din0[176]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  664.775 1.0375 664.91 1.1725 ;
      END
   END din0[176]
   PIN din0[177]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  667.635 1.0375 667.77 1.1725 ;
      END
   END din0[177]
   PIN din0[178]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  670.495 1.0375 670.63 1.1725 ;
      END
   END din0[178]
   PIN din0[179]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  673.355 1.0375 673.49 1.1725 ;
      END
   END din0[179]
   PIN din0[180]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  676.215 1.0375 676.35 1.1725 ;
      END
   END din0[180]
   PIN din0[181]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  679.075 1.0375 679.21 1.1725 ;
      END
   END din0[181]
   PIN din0[182]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  681.935 1.0375 682.07 1.1725 ;
      END
   END din0[182]
   PIN din0[183]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  684.795 1.0375 684.93 1.1725 ;
      END
   END din0[183]
   PIN din0[184]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  687.655 1.0375 687.79 1.1725 ;
      END
   END din0[184]
   PIN din0[185]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  690.515 1.0375 690.65 1.1725 ;
      END
   END din0[185]
   PIN din0[186]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  693.375 1.0375 693.51 1.1725 ;
      END
   END din0[186]
   PIN din0[187]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  696.235 1.0375 696.37 1.1725 ;
      END
   END din0[187]
   PIN din0[188]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  699.095 1.0375 699.23 1.1725 ;
      END
   END din0[188]
   PIN din0[189]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  701.955 1.0375 702.09 1.1725 ;
      END
   END din0[189]
   PIN din0[190]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  704.815 1.0375 704.95 1.1725 ;
      END
   END din0[190]
   PIN din0[191]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  707.675 1.0375 707.81 1.1725 ;
      END
   END din0[191]
   PIN din0[192]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  710.535 1.0375 710.67 1.1725 ;
      END
   END din0[192]
   PIN din0[193]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  713.395 1.0375 713.53 1.1725 ;
      END
   END din0[193]
   PIN din0[194]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  716.255 1.0375 716.39 1.1725 ;
      END
   END din0[194]
   PIN din0[195]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  719.115 1.0375 719.25 1.1725 ;
      END
   END din0[195]
   PIN din0[196]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  721.975 1.0375 722.11 1.1725 ;
      END
   END din0[196]
   PIN din0[197]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  724.835 1.0375 724.97 1.1725 ;
      END
   END din0[197]
   PIN din0[198]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  727.695 1.0375 727.83 1.1725 ;
      END
   END din0[198]
   PIN din0[199]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  730.555 1.0375 730.69 1.1725 ;
      END
   END din0[199]
   PIN din0[200]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  733.415 1.0375 733.55 1.1725 ;
      END
   END din0[200]
   PIN din0[201]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  736.275 1.0375 736.41 1.1725 ;
      END
   END din0[201]
   PIN din0[202]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  739.135 1.0375 739.27 1.1725 ;
      END
   END din0[202]
   PIN din0[203]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  741.995 1.0375 742.13 1.1725 ;
      END
   END din0[203]
   PIN din0[204]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  744.855 1.0375 744.99 1.1725 ;
      END
   END din0[204]
   PIN din0[205]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  747.715 1.0375 747.85 1.1725 ;
      END
   END din0[205]
   PIN din0[206]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  750.575 1.0375 750.71 1.1725 ;
      END
   END din0[206]
   PIN din0[207]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  753.435 1.0375 753.57 1.1725 ;
      END
   END din0[207]
   PIN din0[208]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  756.295 1.0375 756.43 1.1725 ;
      END
   END din0[208]
   PIN din0[209]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  759.155 1.0375 759.29 1.1725 ;
      END
   END din0[209]
   PIN din0[210]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  762.015 1.0375 762.15 1.1725 ;
      END
   END din0[210]
   PIN din0[211]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  764.875 1.0375 765.01 1.1725 ;
      END
   END din0[211]
   PIN din0[212]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  767.735 1.0375 767.87 1.1725 ;
      END
   END din0[212]
   PIN din0[213]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  770.595 1.0375 770.73 1.1725 ;
      END
   END din0[213]
   PIN din0[214]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  773.455 1.0375 773.59 1.1725 ;
      END
   END din0[214]
   PIN din0[215]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  776.315 1.0375 776.45 1.1725 ;
      END
   END din0[215]
   PIN din0[216]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  779.175 1.0375 779.31 1.1725 ;
      END
   END din0[216]
   PIN din0[217]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  782.035 1.0375 782.17 1.1725 ;
      END
   END din0[217]
   PIN din0[218]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  784.895 1.0375 785.03 1.1725 ;
      END
   END din0[218]
   PIN din0[219]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  787.755 1.0375 787.89 1.1725 ;
      END
   END din0[219]
   PIN din0[220]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  790.615 1.0375 790.75 1.1725 ;
      END
   END din0[220]
   PIN din0[221]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  793.475 1.0375 793.61 1.1725 ;
      END
   END din0[221]
   PIN din0[222]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  796.335 1.0375 796.47 1.1725 ;
      END
   END din0[222]
   PIN din0[223]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  799.195 1.0375 799.33 1.1725 ;
      END
   END din0[223]
   PIN din0[224]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  802.055 1.0375 802.19 1.1725 ;
      END
   END din0[224]
   PIN din0[225]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  804.915 1.0375 805.05 1.1725 ;
      END
   END din0[225]
   PIN din0[226]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  807.775 1.0375 807.91 1.1725 ;
      END
   END din0[226]
   PIN din0[227]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  810.635 1.0375 810.77 1.1725 ;
      END
   END din0[227]
   PIN din0[228]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  813.495 1.0375 813.63 1.1725 ;
      END
   END din0[228]
   PIN din0[229]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  816.355 1.0375 816.49 1.1725 ;
      END
   END din0[229]
   PIN din0[230]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  819.215 1.0375 819.35 1.1725 ;
      END
   END din0[230]
   PIN din0[231]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  822.075 1.0375 822.21 1.1725 ;
      END
   END din0[231]
   PIN din0[232]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  824.935 1.0375 825.07 1.1725 ;
      END
   END din0[232]
   PIN din0[233]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  827.795 1.0375 827.93 1.1725 ;
      END
   END din0[233]
   PIN din0[234]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  830.655 1.0375 830.79 1.1725 ;
      END
   END din0[234]
   PIN din0[235]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  833.515 1.0375 833.65 1.1725 ;
      END
   END din0[235]
   PIN din0[236]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  836.375 1.0375 836.51 1.1725 ;
      END
   END din0[236]
   PIN din0[237]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  839.235 1.0375 839.37 1.1725 ;
      END
   END din0[237]
   PIN din0[238]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  842.095 1.0375 842.23 1.1725 ;
      END
   END din0[238]
   PIN din0[239]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  844.955 1.0375 845.09 1.1725 ;
      END
   END din0[239]
   PIN din0[240]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  847.815 1.0375 847.95 1.1725 ;
      END
   END din0[240]
   PIN din0[241]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  850.675 1.0375 850.81 1.1725 ;
      END
   END din0[241]
   PIN din0[242]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  853.535 1.0375 853.67 1.1725 ;
      END
   END din0[242]
   PIN din0[243]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  856.395 1.0375 856.53 1.1725 ;
      END
   END din0[243]
   PIN din0[244]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  859.255 1.0375 859.39 1.1725 ;
      END
   END din0[244]
   PIN din0[245]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  862.115 1.0375 862.25 1.1725 ;
      END
   END din0[245]
   PIN din0[246]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  864.975 1.0375 865.11 1.1725 ;
      END
   END din0[246]
   PIN din0[247]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  867.835 1.0375 867.97 1.1725 ;
      END
   END din0[247]
   PIN din0[248]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  870.695 1.0375 870.83 1.1725 ;
      END
   END din0[248]
   PIN din0[249]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  873.555 1.0375 873.69 1.1725 ;
      END
   END din0[249]
   PIN din0[250]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  876.415 1.0375 876.55 1.1725 ;
      END
   END din0[250]
   PIN din0[251]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  879.275 1.0375 879.41 1.1725 ;
      END
   END din0[251]
   PIN din0[252]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  882.135 1.0375 882.27 1.1725 ;
      END
   END din0[252]
   PIN din0[253]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  884.995 1.0375 885.13 1.1725 ;
      END
   END din0[253]
   PIN din0[254]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  887.855 1.0375 887.99 1.1725 ;
      END
   END din0[254]
   PIN din0[255]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  890.715 1.0375 890.85 1.1725 ;
      END
   END din0[255]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.175 97.17 64.31 97.305 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.175 99.9 64.31 100.035 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.175 102.11 64.31 102.245 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.175 104.84 64.31 104.975 ;
      END
   END addr0[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 60.64 0.42 60.775 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 63.37 0.42 63.505 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.5275 60.725 6.6625 60.86 ;
      END
   END clk0
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.895 1.0375 70.03 1.1725 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.755 1.0375 72.89 1.1725 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.615 1.0375 75.75 1.1725 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.475 1.0375 78.61 1.1725 ;
      END
   END wmask0[3]
   PIN wmask0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.335 1.0375 81.47 1.1725 ;
      END
   END wmask0[4]
   PIN wmask0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  84.195 1.0375 84.33 1.1725 ;
      END
   END wmask0[5]
   PIN wmask0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  87.055 1.0375 87.19 1.1725 ;
      END
   END wmask0[6]
   PIN wmask0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.915 1.0375 90.05 1.1725 ;
      END
   END wmask0[7]
   PIN wmask0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.775 1.0375 92.91 1.1725 ;
      END
   END wmask0[8]
   PIN wmask0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.635 1.0375 95.77 1.1725 ;
      END
   END wmask0[9]
   PIN wmask0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.495 1.0375 98.63 1.1725 ;
      END
   END wmask0[10]
   PIN wmask0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.355 1.0375 101.49 1.1725 ;
      END
   END wmask0[11]
   PIN wmask0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.215 1.0375 104.35 1.1725 ;
      END
   END wmask0[12]
   PIN wmask0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  107.075 1.0375 107.21 1.1725 ;
      END
   END wmask0[13]
   PIN wmask0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.935 1.0375 110.07 1.1725 ;
      END
   END wmask0[14]
   PIN wmask0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  112.795 1.0375 112.93 1.1725 ;
      END
   END wmask0[15]
   PIN wmask0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  115.655 1.0375 115.79 1.1725 ;
      END
   END wmask0[16]
   PIN wmask0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.515 1.0375 118.65 1.1725 ;
      END
   END wmask0[17]
   PIN wmask0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  121.375 1.0375 121.51 1.1725 ;
      END
   END wmask0[18]
   PIN wmask0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  124.235 1.0375 124.37 1.1725 ;
      END
   END wmask0[19]
   PIN wmask0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  127.095 1.0375 127.23 1.1725 ;
      END
   END wmask0[20]
   PIN wmask0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.955 1.0375 130.09 1.1725 ;
      END
   END wmask0[21]
   PIN wmask0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.815 1.0375 132.95 1.1725 ;
      END
   END wmask0[22]
   PIN wmask0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.675 1.0375 135.81 1.1725 ;
      END
   END wmask0[23]
   PIN wmask0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  138.535 1.0375 138.67 1.1725 ;
      END
   END wmask0[24]
   PIN wmask0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  141.395 1.0375 141.53 1.1725 ;
      END
   END wmask0[25]
   PIN wmask0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  144.255 1.0375 144.39 1.1725 ;
      END
   END wmask0[26]
   PIN wmask0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  147.115 1.0375 147.25 1.1725 ;
      END
   END wmask0[27]
   PIN wmask0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.975 1.0375 150.11 1.1725 ;
      END
   END wmask0[28]
   PIN wmask0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.835 1.0375 152.97 1.1725 ;
      END
   END wmask0[29]
   PIN wmask0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  155.695 1.0375 155.83 1.1725 ;
      END
   END wmask0[30]
   PIN wmask0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  158.555 1.0375 158.69 1.1725 ;
      END
   END wmask0[31]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.545 71.7825 92.68 71.9175 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  93.25 71.7825 93.385 71.9175 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  93.955 71.7825 94.09 71.9175 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.66 71.7825 94.795 71.9175 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.365 71.7825 95.5 71.9175 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.07 71.7825 96.205 71.9175 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.775 71.7825 96.91 71.9175 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.48 71.7825 97.615 71.9175 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.185 71.7825 98.32 71.9175 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.89 71.7825 99.025 71.9175 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.595 71.7825 99.73 71.9175 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.3 71.7825 100.435 71.9175 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.005 71.7825 101.14 71.9175 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.71 71.7825 101.845 71.9175 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  102.415 71.7825 102.55 71.9175 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.12 71.7825 103.255 71.9175 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.825 71.7825 103.96 71.9175 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.53 71.7825 104.665 71.9175 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  105.235 71.7825 105.37 71.9175 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  105.94 71.7825 106.075 71.9175 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.645 71.7825 106.78 71.9175 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  107.35 71.7825 107.485 71.9175 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.055 71.7825 108.19 71.9175 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.76 71.7825 108.895 71.9175 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.465 71.7825 109.6 71.9175 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  110.17 71.7825 110.305 71.9175 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  110.875 71.7825 111.01 71.9175 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.58 71.7825 111.715 71.9175 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  112.285 71.7825 112.42 71.9175 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  112.99 71.7825 113.125 71.9175 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.695 71.7825 113.83 71.9175 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.4 71.7825 114.535 71.9175 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  115.105 71.7825 115.24 71.9175 ;
      END
   END dout0[32]
   PIN dout0[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  115.81 71.7825 115.945 71.9175 ;
      END
   END dout0[33]
   PIN dout0[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  116.515 71.7825 116.65 71.9175 ;
      END
   END dout0[34]
   PIN dout0[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  117.22 71.7825 117.355 71.9175 ;
      END
   END dout0[35]
   PIN dout0[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  117.925 71.7825 118.06 71.9175 ;
      END
   END dout0[36]
   PIN dout0[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.63 71.7825 118.765 71.9175 ;
      END
   END dout0[37]
   PIN dout0[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  119.335 71.7825 119.47 71.9175 ;
      END
   END dout0[38]
   PIN dout0[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.04 71.7825 120.175 71.9175 ;
      END
   END dout0[39]
   PIN dout0[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.745 71.7825 120.88 71.9175 ;
      END
   END dout0[40]
   PIN dout0[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  121.45 71.7825 121.585 71.9175 ;
      END
   END dout0[41]
   PIN dout0[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  122.155 71.7825 122.29 71.9175 ;
      END
   END dout0[42]
   PIN dout0[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  122.86 71.7825 122.995 71.9175 ;
      END
   END dout0[43]
   PIN dout0[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.565 71.7825 123.7 71.9175 ;
      END
   END dout0[44]
   PIN dout0[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  124.27 71.7825 124.405 71.9175 ;
      END
   END dout0[45]
   PIN dout0[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  124.975 71.7825 125.11 71.9175 ;
      END
   END dout0[46]
   PIN dout0[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  125.68 71.7825 125.815 71.9175 ;
      END
   END dout0[47]
   PIN dout0[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.385 71.7825 126.52 71.9175 ;
      END
   END dout0[48]
   PIN dout0[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  127.09 71.7825 127.225 71.9175 ;
      END
   END dout0[49]
   PIN dout0[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  127.795 71.7825 127.93 71.9175 ;
      END
   END dout0[50]
   PIN dout0[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  128.5 71.7825 128.635 71.9175 ;
      END
   END dout0[51]
   PIN dout0[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.205 71.7825 129.34 71.9175 ;
      END
   END dout0[52]
   PIN dout0[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.91 71.7825 130.045 71.9175 ;
      END
   END dout0[53]
   PIN dout0[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  130.615 71.7825 130.75 71.9175 ;
      END
   END dout0[54]
   PIN dout0[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.32 71.7825 131.455 71.9175 ;
      END
   END dout0[55]
   PIN dout0[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.025 71.7825 132.16 71.9175 ;
      END
   END dout0[56]
   PIN dout0[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.73 71.7825 132.865 71.9175 ;
      END
   END dout0[57]
   PIN dout0[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  133.435 71.7825 133.57 71.9175 ;
      END
   END dout0[58]
   PIN dout0[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.14 71.7825 134.275 71.9175 ;
      END
   END dout0[59]
   PIN dout0[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.845 71.7825 134.98 71.9175 ;
      END
   END dout0[60]
   PIN dout0[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.55 71.7825 135.685 71.9175 ;
      END
   END dout0[61]
   PIN dout0[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  136.255 71.7825 136.39 71.9175 ;
      END
   END dout0[62]
   PIN dout0[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  136.96 71.7825 137.095 71.9175 ;
      END
   END dout0[63]
   PIN dout0[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.665 71.7825 137.8 71.9175 ;
      END
   END dout0[64]
   PIN dout0[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  138.37 71.7825 138.505 71.9175 ;
      END
   END dout0[65]
   PIN dout0[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  139.075 71.7825 139.21 71.9175 ;
      END
   END dout0[66]
   PIN dout0[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  139.78 71.7825 139.915 71.9175 ;
      END
   END dout0[67]
   PIN dout0[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.485 71.7825 140.62 71.9175 ;
      END
   END dout0[68]
   PIN dout0[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  141.19 71.7825 141.325 71.9175 ;
      END
   END dout0[69]
   PIN dout0[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  141.895 71.7825 142.03 71.9175 ;
      END
   END dout0[70]
   PIN dout0[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  142.6 71.7825 142.735 71.9175 ;
      END
   END dout0[71]
   PIN dout0[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.305 71.7825 143.44 71.9175 ;
      END
   END dout0[72]
   PIN dout0[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  144.01 71.7825 144.145 71.9175 ;
      END
   END dout0[73]
   PIN dout0[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  144.715 71.7825 144.85 71.9175 ;
      END
   END dout0[74]
   PIN dout0[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  145.42 71.7825 145.555 71.9175 ;
      END
   END dout0[75]
   PIN dout0[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.125 71.7825 146.26 71.9175 ;
      END
   END dout0[76]
   PIN dout0[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.83 71.7825 146.965 71.9175 ;
      END
   END dout0[77]
   PIN dout0[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  147.535 71.7825 147.67 71.9175 ;
      END
   END dout0[78]
   PIN dout0[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  148.24 71.7825 148.375 71.9175 ;
      END
   END dout0[79]
   PIN dout0[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  148.945 71.7825 149.08 71.9175 ;
      END
   END dout0[80]
   PIN dout0[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.65 71.7825 149.785 71.9175 ;
      END
   END dout0[81]
   PIN dout0[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  150.355 71.7825 150.49 71.9175 ;
      END
   END dout0[82]
   PIN dout0[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  151.06 71.7825 151.195 71.9175 ;
      END
   END dout0[83]
   PIN dout0[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  151.765 71.7825 151.9 71.9175 ;
      END
   END dout0[84]
   PIN dout0[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  152.47 71.7825 152.605 71.9175 ;
      END
   END dout0[85]
   PIN dout0[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  153.175 71.7825 153.31 71.9175 ;
      END
   END dout0[86]
   PIN dout0[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  153.88 71.7825 154.015 71.9175 ;
      END
   END dout0[87]
   PIN dout0[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.585 71.7825 154.72 71.9175 ;
      END
   END dout0[88]
   PIN dout0[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  155.29 71.7825 155.425 71.9175 ;
      END
   END dout0[89]
   PIN dout0[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  155.995 71.7825 156.13 71.9175 ;
      END
   END dout0[90]
   PIN dout0[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  156.7 71.7825 156.835 71.9175 ;
      END
   END dout0[91]
   PIN dout0[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  157.405 71.7825 157.54 71.9175 ;
      END
   END dout0[92]
   PIN dout0[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  158.11 71.7825 158.245 71.9175 ;
      END
   END dout0[93]
   PIN dout0[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  158.815 71.7825 158.95 71.9175 ;
      END
   END dout0[94]
   PIN dout0[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  159.52 71.7825 159.655 71.9175 ;
      END
   END dout0[95]
   PIN dout0[96]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.225 71.7825 160.36 71.9175 ;
      END
   END dout0[96]
   PIN dout0[97]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.93 71.7825 161.065 71.9175 ;
      END
   END dout0[97]
   PIN dout0[98]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  161.635 71.7825 161.77 71.9175 ;
      END
   END dout0[98]
   PIN dout0[99]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  162.34 71.7825 162.475 71.9175 ;
      END
   END dout0[99]
   PIN dout0[100]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.045 71.7825 163.18 71.9175 ;
      END
   END dout0[100]
   PIN dout0[101]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.75 71.7825 163.885 71.9175 ;
      END
   END dout0[101]
   PIN dout0[102]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  164.455 71.7825 164.59 71.9175 ;
      END
   END dout0[102]
   PIN dout0[103]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  165.16 71.7825 165.295 71.9175 ;
      END
   END dout0[103]
   PIN dout0[104]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  165.865 71.7825 166.0 71.9175 ;
      END
   END dout0[104]
   PIN dout0[105]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.57 71.7825 166.705 71.9175 ;
      END
   END dout0[105]
   PIN dout0[106]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  167.275 71.7825 167.41 71.9175 ;
      END
   END dout0[106]
   PIN dout0[107]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  167.98 71.7825 168.115 71.9175 ;
      END
   END dout0[107]
   PIN dout0[108]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  168.685 71.7825 168.82 71.9175 ;
      END
   END dout0[108]
   PIN dout0[109]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.39 71.7825 169.525 71.9175 ;
      END
   END dout0[109]
   PIN dout0[110]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  170.095 71.7825 170.23 71.9175 ;
      END
   END dout0[110]
   PIN dout0[111]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  170.8 71.7825 170.935 71.9175 ;
      END
   END dout0[111]
   PIN dout0[112]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  171.505 71.7825 171.64 71.9175 ;
      END
   END dout0[112]
   PIN dout0[113]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.21 71.7825 172.345 71.9175 ;
      END
   END dout0[113]
   PIN dout0[114]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  172.915 71.7825 173.05 71.9175 ;
      END
   END dout0[114]
   PIN dout0[115]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  173.62 71.7825 173.755 71.9175 ;
      END
   END dout0[115]
   PIN dout0[116]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.325 71.7825 174.46 71.9175 ;
      END
   END dout0[116]
   PIN dout0[117]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  175.03 71.7825 175.165 71.9175 ;
      END
   END dout0[117]
   PIN dout0[118]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  175.735 71.7825 175.87 71.9175 ;
      END
   END dout0[118]
   PIN dout0[119]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  176.44 71.7825 176.575 71.9175 ;
      END
   END dout0[119]
   PIN dout0[120]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.145 71.7825 177.28 71.9175 ;
      END
   END dout0[120]
   PIN dout0[121]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.85 71.7825 177.985 71.9175 ;
      END
   END dout0[121]
   PIN dout0[122]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  178.555 71.7825 178.69 71.9175 ;
      END
   END dout0[122]
   PIN dout0[123]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.26 71.7825 179.395 71.9175 ;
      END
   END dout0[123]
   PIN dout0[124]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  179.965 71.7825 180.1 71.9175 ;
      END
   END dout0[124]
   PIN dout0[125]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.67 71.7825 180.805 71.9175 ;
      END
   END dout0[125]
   PIN dout0[126]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  181.375 71.7825 181.51 71.9175 ;
      END
   END dout0[126]
   PIN dout0[127]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  182.08 71.7825 182.215 71.9175 ;
      END
   END dout0[127]
   PIN dout0[128]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  182.785 71.7825 182.92 71.9175 ;
      END
   END dout0[128]
   PIN dout0[129]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.49 71.7825 183.625 71.9175 ;
      END
   END dout0[129]
   PIN dout0[130]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  184.195 71.7825 184.33 71.9175 ;
      END
   END dout0[130]
   PIN dout0[131]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  184.9 71.7825 185.035 71.9175 ;
      END
   END dout0[131]
   PIN dout0[132]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  185.605 71.7825 185.74 71.9175 ;
      END
   END dout0[132]
   PIN dout0[133]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.31 71.7825 186.445 71.9175 ;
      END
   END dout0[133]
   PIN dout0[134]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  187.015 71.7825 187.15 71.9175 ;
      END
   END dout0[134]
   PIN dout0[135]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  187.72 71.7825 187.855 71.9175 ;
      END
   END dout0[135]
   PIN dout0[136]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  188.425 71.7825 188.56 71.9175 ;
      END
   END dout0[136]
   PIN dout0[137]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.13 71.7825 189.265 71.9175 ;
      END
   END dout0[137]
   PIN dout0[138]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.835 71.7825 189.97 71.9175 ;
      END
   END dout0[138]
   PIN dout0[139]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  190.54 71.7825 190.675 71.9175 ;
      END
   END dout0[139]
   PIN dout0[140]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  191.245 71.7825 191.38 71.9175 ;
      END
   END dout0[140]
   PIN dout0[141]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  191.95 71.7825 192.085 71.9175 ;
      END
   END dout0[141]
   PIN dout0[142]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  192.655 71.7825 192.79 71.9175 ;
      END
   END dout0[142]
   PIN dout0[143]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  193.36 71.7825 193.495 71.9175 ;
      END
   END dout0[143]
   PIN dout0[144]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  194.065 71.7825 194.2 71.9175 ;
      END
   END dout0[144]
   PIN dout0[145]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  194.77 71.7825 194.905 71.9175 ;
      END
   END dout0[145]
   PIN dout0[146]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  195.475 71.7825 195.61 71.9175 ;
      END
   END dout0[146]
   PIN dout0[147]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  196.18 71.7825 196.315 71.9175 ;
      END
   END dout0[147]
   PIN dout0[148]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  196.885 71.7825 197.02 71.9175 ;
      END
   END dout0[148]
   PIN dout0[149]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  197.59 71.7825 197.725 71.9175 ;
      END
   END dout0[149]
   PIN dout0[150]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  198.295 71.7825 198.43 71.9175 ;
      END
   END dout0[150]
   PIN dout0[151]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  199.0 71.7825 199.135 71.9175 ;
      END
   END dout0[151]
   PIN dout0[152]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  199.705 71.7825 199.84 71.9175 ;
      END
   END dout0[152]
   PIN dout0[153]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  200.41 71.7825 200.545 71.9175 ;
      END
   END dout0[153]
   PIN dout0[154]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  201.115 71.7825 201.25 71.9175 ;
      END
   END dout0[154]
   PIN dout0[155]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  201.82 71.7825 201.955 71.9175 ;
      END
   END dout0[155]
   PIN dout0[156]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  202.525 71.7825 202.66 71.9175 ;
      END
   END dout0[156]
   PIN dout0[157]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  203.23 71.7825 203.365 71.9175 ;
      END
   END dout0[157]
   PIN dout0[158]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  203.935 71.7825 204.07 71.9175 ;
      END
   END dout0[158]
   PIN dout0[159]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  204.64 71.7825 204.775 71.9175 ;
      END
   END dout0[159]
   PIN dout0[160]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  205.345 71.7825 205.48 71.9175 ;
      END
   END dout0[160]
   PIN dout0[161]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  206.05 71.7825 206.185 71.9175 ;
      END
   END dout0[161]
   PIN dout0[162]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  206.755 71.7825 206.89 71.9175 ;
      END
   END dout0[162]
   PIN dout0[163]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  207.46 71.7825 207.595 71.9175 ;
      END
   END dout0[163]
   PIN dout0[164]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  208.165 71.7825 208.3 71.9175 ;
      END
   END dout0[164]
   PIN dout0[165]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  208.87 71.7825 209.005 71.9175 ;
      END
   END dout0[165]
   PIN dout0[166]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  209.575 71.7825 209.71 71.9175 ;
      END
   END dout0[166]
   PIN dout0[167]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  210.28 71.7825 210.415 71.9175 ;
      END
   END dout0[167]
   PIN dout0[168]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  210.985 71.7825 211.12 71.9175 ;
      END
   END dout0[168]
   PIN dout0[169]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  211.69 71.7825 211.825 71.9175 ;
      END
   END dout0[169]
   PIN dout0[170]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  212.395 71.7825 212.53 71.9175 ;
      END
   END dout0[170]
   PIN dout0[171]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  213.1 71.7825 213.235 71.9175 ;
      END
   END dout0[171]
   PIN dout0[172]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  213.805 71.7825 213.94 71.9175 ;
      END
   END dout0[172]
   PIN dout0[173]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  214.51 71.7825 214.645 71.9175 ;
      END
   END dout0[173]
   PIN dout0[174]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  215.215 71.7825 215.35 71.9175 ;
      END
   END dout0[174]
   PIN dout0[175]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  215.92 71.7825 216.055 71.9175 ;
      END
   END dout0[175]
   PIN dout0[176]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  216.625 71.7825 216.76 71.9175 ;
      END
   END dout0[176]
   PIN dout0[177]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  217.33 71.7825 217.465 71.9175 ;
      END
   END dout0[177]
   PIN dout0[178]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  218.035 71.7825 218.17 71.9175 ;
      END
   END dout0[178]
   PIN dout0[179]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  218.74 71.7825 218.875 71.9175 ;
      END
   END dout0[179]
   PIN dout0[180]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  219.445 71.7825 219.58 71.9175 ;
      END
   END dout0[180]
   PIN dout0[181]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  220.15 71.7825 220.285 71.9175 ;
      END
   END dout0[181]
   PIN dout0[182]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  220.855 71.7825 220.99 71.9175 ;
      END
   END dout0[182]
   PIN dout0[183]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  221.56 71.7825 221.695 71.9175 ;
      END
   END dout0[183]
   PIN dout0[184]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  222.265 71.7825 222.4 71.9175 ;
      END
   END dout0[184]
   PIN dout0[185]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  222.97 71.7825 223.105 71.9175 ;
      END
   END dout0[185]
   PIN dout0[186]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  223.675 71.7825 223.81 71.9175 ;
      END
   END dout0[186]
   PIN dout0[187]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  224.38 71.7825 224.515 71.9175 ;
      END
   END dout0[187]
   PIN dout0[188]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  225.085 71.7825 225.22 71.9175 ;
      END
   END dout0[188]
   PIN dout0[189]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  225.79 71.7825 225.925 71.9175 ;
      END
   END dout0[189]
   PIN dout0[190]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  226.495 71.7825 226.63 71.9175 ;
      END
   END dout0[190]
   PIN dout0[191]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  227.2 71.7825 227.335 71.9175 ;
      END
   END dout0[191]
   PIN dout0[192]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  227.905 71.7825 228.04 71.9175 ;
      END
   END dout0[192]
   PIN dout0[193]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  228.61 71.7825 228.745 71.9175 ;
      END
   END dout0[193]
   PIN dout0[194]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  229.315 71.7825 229.45 71.9175 ;
      END
   END dout0[194]
   PIN dout0[195]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  230.02 71.7825 230.155 71.9175 ;
      END
   END dout0[195]
   PIN dout0[196]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  230.725 71.7825 230.86 71.9175 ;
      END
   END dout0[196]
   PIN dout0[197]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  231.43 71.7825 231.565 71.9175 ;
      END
   END dout0[197]
   PIN dout0[198]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  232.135 71.7825 232.27 71.9175 ;
      END
   END dout0[198]
   PIN dout0[199]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  232.84 71.7825 232.975 71.9175 ;
      END
   END dout0[199]
   PIN dout0[200]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  233.545 71.7825 233.68 71.9175 ;
      END
   END dout0[200]
   PIN dout0[201]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  234.25 71.7825 234.385 71.9175 ;
      END
   END dout0[201]
   PIN dout0[202]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  234.955 71.7825 235.09 71.9175 ;
      END
   END dout0[202]
   PIN dout0[203]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  235.66 71.7825 235.795 71.9175 ;
      END
   END dout0[203]
   PIN dout0[204]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  236.365 71.7825 236.5 71.9175 ;
      END
   END dout0[204]
   PIN dout0[205]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  237.07 71.7825 237.205 71.9175 ;
      END
   END dout0[205]
   PIN dout0[206]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  237.775 71.7825 237.91 71.9175 ;
      END
   END dout0[206]
   PIN dout0[207]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  238.48 71.7825 238.615 71.9175 ;
      END
   END dout0[207]
   PIN dout0[208]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  239.185 71.7825 239.32 71.9175 ;
      END
   END dout0[208]
   PIN dout0[209]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  239.89 71.7825 240.025 71.9175 ;
      END
   END dout0[209]
   PIN dout0[210]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  240.595 71.7825 240.73 71.9175 ;
      END
   END dout0[210]
   PIN dout0[211]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  241.3 71.7825 241.435 71.9175 ;
      END
   END dout0[211]
   PIN dout0[212]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  242.005 71.7825 242.14 71.9175 ;
      END
   END dout0[212]
   PIN dout0[213]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  242.71 71.7825 242.845 71.9175 ;
      END
   END dout0[213]
   PIN dout0[214]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  243.415 71.7825 243.55 71.9175 ;
      END
   END dout0[214]
   PIN dout0[215]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  244.12 71.7825 244.255 71.9175 ;
      END
   END dout0[215]
   PIN dout0[216]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  244.825 71.7825 244.96 71.9175 ;
      END
   END dout0[216]
   PIN dout0[217]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  245.53 71.7825 245.665 71.9175 ;
      END
   END dout0[217]
   PIN dout0[218]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  246.235 71.7825 246.37 71.9175 ;
      END
   END dout0[218]
   PIN dout0[219]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  246.94 71.7825 247.075 71.9175 ;
      END
   END dout0[219]
   PIN dout0[220]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  247.645 71.7825 247.78 71.9175 ;
      END
   END dout0[220]
   PIN dout0[221]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  248.35 71.7825 248.485 71.9175 ;
      END
   END dout0[221]
   PIN dout0[222]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  249.055 71.7825 249.19 71.9175 ;
      END
   END dout0[222]
   PIN dout0[223]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  249.76 71.7825 249.895 71.9175 ;
      END
   END dout0[223]
   PIN dout0[224]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  250.465 71.7825 250.6 71.9175 ;
      END
   END dout0[224]
   PIN dout0[225]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  251.17 71.7825 251.305 71.9175 ;
      END
   END dout0[225]
   PIN dout0[226]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  251.875 71.7825 252.01 71.9175 ;
      END
   END dout0[226]
   PIN dout0[227]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  252.58 71.7825 252.715 71.9175 ;
      END
   END dout0[227]
   PIN dout0[228]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  253.285 71.7825 253.42 71.9175 ;
      END
   END dout0[228]
   PIN dout0[229]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  253.99 71.7825 254.125 71.9175 ;
      END
   END dout0[229]
   PIN dout0[230]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  254.695 71.7825 254.83 71.9175 ;
      END
   END dout0[230]
   PIN dout0[231]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  255.4 71.7825 255.535 71.9175 ;
      END
   END dout0[231]
   PIN dout0[232]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  256.105 71.7825 256.24 71.9175 ;
      END
   END dout0[232]
   PIN dout0[233]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  256.81 71.7825 256.945 71.9175 ;
      END
   END dout0[233]
   PIN dout0[234]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  257.515 71.7825 257.65 71.9175 ;
      END
   END dout0[234]
   PIN dout0[235]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  258.22 71.7825 258.355 71.9175 ;
      END
   END dout0[235]
   PIN dout0[236]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  258.925 71.7825 259.06 71.9175 ;
      END
   END dout0[236]
   PIN dout0[237]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  259.63 71.7825 259.765 71.9175 ;
      END
   END dout0[237]
   PIN dout0[238]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  260.335 71.7825 260.47 71.9175 ;
      END
   END dout0[238]
   PIN dout0[239]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  261.04 71.7825 261.175 71.9175 ;
      END
   END dout0[239]
   PIN dout0[240]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  261.745 71.7825 261.88 71.9175 ;
      END
   END dout0[240]
   PIN dout0[241]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  262.45 71.7825 262.585 71.9175 ;
      END
   END dout0[241]
   PIN dout0[242]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  263.155 71.7825 263.29 71.9175 ;
      END
   END dout0[242]
   PIN dout0[243]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  263.86 71.7825 263.995 71.9175 ;
      END
   END dout0[243]
   PIN dout0[244]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  264.565 71.7825 264.7 71.9175 ;
      END
   END dout0[244]
   PIN dout0[245]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  265.27 71.7825 265.405 71.9175 ;
      END
   END dout0[245]
   PIN dout0[246]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  265.975 71.7825 266.11 71.9175 ;
      END
   END dout0[246]
   PIN dout0[247]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  266.68 71.7825 266.815 71.9175 ;
      END
   END dout0[247]
   PIN dout0[248]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  267.385 71.7825 267.52 71.9175 ;
      END
   END dout0[248]
   PIN dout0[249]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  268.09 71.7825 268.225 71.9175 ;
      END
   END dout0[249]
   PIN dout0[250]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  268.795 71.7825 268.93 71.9175 ;
      END
   END dout0[250]
   PIN dout0[251]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  269.5 71.7825 269.635 71.9175 ;
      END
   END dout0[251]
   PIN dout0[252]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  270.205 71.7825 270.34 71.9175 ;
      END
   END dout0[252]
   PIN dout0[253]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  270.91 71.7825 271.045 71.9175 ;
      END
   END dout0[253]
   PIN dout0[254]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  271.615 71.7825 271.75 71.9175 ;
      END
   END dout0[254]
   PIN dout0[255]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  272.32 71.7825 272.455 71.9175 ;
      END
   END dout0[255]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 893.22 124.97 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 893.22 124.97 ;
   LAYER  metal3 ;
      RECT  0.14 0.14 161.275 0.8975 ;
      RECT  161.275 0.14 161.69 0.8975 ;
      RECT  161.69 0.14 893.22 0.8975 ;
      RECT  161.69 0.8975 164.135 1.3125 ;
      RECT  164.55 0.8975 166.995 1.3125 ;
      RECT  167.41 0.8975 169.855 1.3125 ;
      RECT  170.27 0.8975 172.715 1.3125 ;
      RECT  173.13 0.8975 175.575 1.3125 ;
      RECT  175.99 0.8975 178.435 1.3125 ;
      RECT  178.85 0.8975 181.295 1.3125 ;
      RECT  181.71 0.8975 184.155 1.3125 ;
      RECT  184.57 0.8975 187.015 1.3125 ;
      RECT  187.43 0.8975 189.875 1.3125 ;
      RECT  190.29 0.8975 192.735 1.3125 ;
      RECT  193.15 0.8975 195.595 1.3125 ;
      RECT  196.01 0.8975 198.455 1.3125 ;
      RECT  198.87 0.8975 201.315 1.3125 ;
      RECT  201.73 0.8975 204.175 1.3125 ;
      RECT  204.59 0.8975 207.035 1.3125 ;
      RECT  207.45 0.8975 209.895 1.3125 ;
      RECT  210.31 0.8975 212.755 1.3125 ;
      RECT  213.17 0.8975 215.615 1.3125 ;
      RECT  216.03 0.8975 218.475 1.3125 ;
      RECT  218.89 0.8975 221.335 1.3125 ;
      RECT  221.75 0.8975 224.195 1.3125 ;
      RECT  224.61 0.8975 227.055 1.3125 ;
      RECT  227.47 0.8975 229.915 1.3125 ;
      RECT  230.33 0.8975 232.775 1.3125 ;
      RECT  233.19 0.8975 235.635 1.3125 ;
      RECT  236.05 0.8975 238.495 1.3125 ;
      RECT  238.91 0.8975 241.355 1.3125 ;
      RECT  241.77 0.8975 244.215 1.3125 ;
      RECT  244.63 0.8975 247.075 1.3125 ;
      RECT  247.49 0.8975 249.935 1.3125 ;
      RECT  250.35 0.8975 252.795 1.3125 ;
      RECT  253.21 0.8975 255.655 1.3125 ;
      RECT  256.07 0.8975 258.515 1.3125 ;
      RECT  258.93 0.8975 261.375 1.3125 ;
      RECT  261.79 0.8975 264.235 1.3125 ;
      RECT  264.65 0.8975 267.095 1.3125 ;
      RECT  267.51 0.8975 269.955 1.3125 ;
      RECT  270.37 0.8975 272.815 1.3125 ;
      RECT  273.23 0.8975 275.675 1.3125 ;
      RECT  276.09 0.8975 278.535 1.3125 ;
      RECT  278.95 0.8975 281.395 1.3125 ;
      RECT  281.81 0.8975 284.255 1.3125 ;
      RECT  284.67 0.8975 287.115 1.3125 ;
      RECT  287.53 0.8975 289.975 1.3125 ;
      RECT  290.39 0.8975 292.835 1.3125 ;
      RECT  293.25 0.8975 295.695 1.3125 ;
      RECT  296.11 0.8975 298.555 1.3125 ;
      RECT  298.97 0.8975 301.415 1.3125 ;
      RECT  301.83 0.8975 304.275 1.3125 ;
      RECT  304.69 0.8975 307.135 1.3125 ;
      RECT  307.55 0.8975 309.995 1.3125 ;
      RECT  310.41 0.8975 312.855 1.3125 ;
      RECT  313.27 0.8975 315.715 1.3125 ;
      RECT  316.13 0.8975 318.575 1.3125 ;
      RECT  318.99 0.8975 321.435 1.3125 ;
      RECT  321.85 0.8975 324.295 1.3125 ;
      RECT  324.71 0.8975 327.155 1.3125 ;
      RECT  327.57 0.8975 330.015 1.3125 ;
      RECT  330.43 0.8975 332.875 1.3125 ;
      RECT  333.29 0.8975 335.735 1.3125 ;
      RECT  336.15 0.8975 338.595 1.3125 ;
      RECT  339.01 0.8975 341.455 1.3125 ;
      RECT  341.87 0.8975 344.315 1.3125 ;
      RECT  344.73 0.8975 347.175 1.3125 ;
      RECT  347.59 0.8975 350.035 1.3125 ;
      RECT  350.45 0.8975 352.895 1.3125 ;
      RECT  353.31 0.8975 355.755 1.3125 ;
      RECT  356.17 0.8975 358.615 1.3125 ;
      RECT  359.03 0.8975 361.475 1.3125 ;
      RECT  361.89 0.8975 364.335 1.3125 ;
      RECT  364.75 0.8975 367.195 1.3125 ;
      RECT  367.61 0.8975 370.055 1.3125 ;
      RECT  370.47 0.8975 372.915 1.3125 ;
      RECT  373.33 0.8975 375.775 1.3125 ;
      RECT  376.19 0.8975 378.635 1.3125 ;
      RECT  379.05 0.8975 381.495 1.3125 ;
      RECT  381.91 0.8975 384.355 1.3125 ;
      RECT  384.77 0.8975 387.215 1.3125 ;
      RECT  387.63 0.8975 390.075 1.3125 ;
      RECT  390.49 0.8975 392.935 1.3125 ;
      RECT  393.35 0.8975 395.795 1.3125 ;
      RECT  396.21 0.8975 398.655 1.3125 ;
      RECT  399.07 0.8975 401.515 1.3125 ;
      RECT  401.93 0.8975 404.375 1.3125 ;
      RECT  404.79 0.8975 407.235 1.3125 ;
      RECT  407.65 0.8975 410.095 1.3125 ;
      RECT  410.51 0.8975 412.955 1.3125 ;
      RECT  413.37 0.8975 415.815 1.3125 ;
      RECT  416.23 0.8975 418.675 1.3125 ;
      RECT  419.09 0.8975 421.535 1.3125 ;
      RECT  421.95 0.8975 424.395 1.3125 ;
      RECT  424.81 0.8975 427.255 1.3125 ;
      RECT  427.67 0.8975 430.115 1.3125 ;
      RECT  430.53 0.8975 432.975 1.3125 ;
      RECT  433.39 0.8975 435.835 1.3125 ;
      RECT  436.25 0.8975 438.695 1.3125 ;
      RECT  439.11 0.8975 441.555 1.3125 ;
      RECT  441.97 0.8975 444.415 1.3125 ;
      RECT  444.83 0.8975 447.275 1.3125 ;
      RECT  447.69 0.8975 450.135 1.3125 ;
      RECT  450.55 0.8975 452.995 1.3125 ;
      RECT  453.41 0.8975 455.855 1.3125 ;
      RECT  456.27 0.8975 458.715 1.3125 ;
      RECT  459.13 0.8975 461.575 1.3125 ;
      RECT  461.99 0.8975 464.435 1.3125 ;
      RECT  464.85 0.8975 467.295 1.3125 ;
      RECT  467.71 0.8975 470.155 1.3125 ;
      RECT  470.57 0.8975 473.015 1.3125 ;
      RECT  473.43 0.8975 475.875 1.3125 ;
      RECT  476.29 0.8975 478.735 1.3125 ;
      RECT  479.15 0.8975 481.595 1.3125 ;
      RECT  482.01 0.8975 484.455 1.3125 ;
      RECT  484.87 0.8975 487.315 1.3125 ;
      RECT  487.73 0.8975 490.175 1.3125 ;
      RECT  490.59 0.8975 493.035 1.3125 ;
      RECT  493.45 0.8975 495.895 1.3125 ;
      RECT  496.31 0.8975 498.755 1.3125 ;
      RECT  499.17 0.8975 501.615 1.3125 ;
      RECT  502.03 0.8975 504.475 1.3125 ;
      RECT  504.89 0.8975 507.335 1.3125 ;
      RECT  507.75 0.8975 510.195 1.3125 ;
      RECT  510.61 0.8975 513.055 1.3125 ;
      RECT  513.47 0.8975 515.915 1.3125 ;
      RECT  516.33 0.8975 518.775 1.3125 ;
      RECT  519.19 0.8975 521.635 1.3125 ;
      RECT  522.05 0.8975 524.495 1.3125 ;
      RECT  524.91 0.8975 527.355 1.3125 ;
      RECT  527.77 0.8975 530.215 1.3125 ;
      RECT  530.63 0.8975 533.075 1.3125 ;
      RECT  533.49 0.8975 535.935 1.3125 ;
      RECT  536.35 0.8975 538.795 1.3125 ;
      RECT  539.21 0.8975 541.655 1.3125 ;
      RECT  542.07 0.8975 544.515 1.3125 ;
      RECT  544.93 0.8975 547.375 1.3125 ;
      RECT  547.79 0.8975 550.235 1.3125 ;
      RECT  550.65 0.8975 553.095 1.3125 ;
      RECT  553.51 0.8975 555.955 1.3125 ;
      RECT  556.37 0.8975 558.815 1.3125 ;
      RECT  559.23 0.8975 561.675 1.3125 ;
      RECT  562.09 0.8975 564.535 1.3125 ;
      RECT  564.95 0.8975 567.395 1.3125 ;
      RECT  567.81 0.8975 570.255 1.3125 ;
      RECT  570.67 0.8975 573.115 1.3125 ;
      RECT  573.53 0.8975 575.975 1.3125 ;
      RECT  576.39 0.8975 578.835 1.3125 ;
      RECT  579.25 0.8975 581.695 1.3125 ;
      RECT  582.11 0.8975 584.555 1.3125 ;
      RECT  584.97 0.8975 587.415 1.3125 ;
      RECT  587.83 0.8975 590.275 1.3125 ;
      RECT  590.69 0.8975 593.135 1.3125 ;
      RECT  593.55 0.8975 595.995 1.3125 ;
      RECT  596.41 0.8975 598.855 1.3125 ;
      RECT  599.27 0.8975 601.715 1.3125 ;
      RECT  602.13 0.8975 604.575 1.3125 ;
      RECT  604.99 0.8975 607.435 1.3125 ;
      RECT  607.85 0.8975 610.295 1.3125 ;
      RECT  610.71 0.8975 613.155 1.3125 ;
      RECT  613.57 0.8975 616.015 1.3125 ;
      RECT  616.43 0.8975 618.875 1.3125 ;
      RECT  619.29 0.8975 621.735 1.3125 ;
      RECT  622.15 0.8975 624.595 1.3125 ;
      RECT  625.01 0.8975 627.455 1.3125 ;
      RECT  627.87 0.8975 630.315 1.3125 ;
      RECT  630.73 0.8975 633.175 1.3125 ;
      RECT  633.59 0.8975 636.035 1.3125 ;
      RECT  636.45 0.8975 638.895 1.3125 ;
      RECT  639.31 0.8975 641.755 1.3125 ;
      RECT  642.17 0.8975 644.615 1.3125 ;
      RECT  645.03 0.8975 647.475 1.3125 ;
      RECT  647.89 0.8975 650.335 1.3125 ;
      RECT  650.75 0.8975 653.195 1.3125 ;
      RECT  653.61 0.8975 656.055 1.3125 ;
      RECT  656.47 0.8975 658.915 1.3125 ;
      RECT  659.33 0.8975 661.775 1.3125 ;
      RECT  662.19 0.8975 664.635 1.3125 ;
      RECT  665.05 0.8975 667.495 1.3125 ;
      RECT  667.91 0.8975 670.355 1.3125 ;
      RECT  670.77 0.8975 673.215 1.3125 ;
      RECT  673.63 0.8975 676.075 1.3125 ;
      RECT  676.49 0.8975 678.935 1.3125 ;
      RECT  679.35 0.8975 681.795 1.3125 ;
      RECT  682.21 0.8975 684.655 1.3125 ;
      RECT  685.07 0.8975 687.515 1.3125 ;
      RECT  687.93 0.8975 690.375 1.3125 ;
      RECT  690.79 0.8975 693.235 1.3125 ;
      RECT  693.65 0.8975 696.095 1.3125 ;
      RECT  696.51 0.8975 698.955 1.3125 ;
      RECT  699.37 0.8975 701.815 1.3125 ;
      RECT  702.23 0.8975 704.675 1.3125 ;
      RECT  705.09 0.8975 707.535 1.3125 ;
      RECT  707.95 0.8975 710.395 1.3125 ;
      RECT  710.81 0.8975 713.255 1.3125 ;
      RECT  713.67 0.8975 716.115 1.3125 ;
      RECT  716.53 0.8975 718.975 1.3125 ;
      RECT  719.39 0.8975 721.835 1.3125 ;
      RECT  722.25 0.8975 724.695 1.3125 ;
      RECT  725.11 0.8975 727.555 1.3125 ;
      RECT  727.97 0.8975 730.415 1.3125 ;
      RECT  730.83 0.8975 733.275 1.3125 ;
      RECT  733.69 0.8975 736.135 1.3125 ;
      RECT  736.55 0.8975 738.995 1.3125 ;
      RECT  739.41 0.8975 741.855 1.3125 ;
      RECT  742.27 0.8975 744.715 1.3125 ;
      RECT  745.13 0.8975 747.575 1.3125 ;
      RECT  747.99 0.8975 750.435 1.3125 ;
      RECT  750.85 0.8975 753.295 1.3125 ;
      RECT  753.71 0.8975 756.155 1.3125 ;
      RECT  756.57 0.8975 759.015 1.3125 ;
      RECT  759.43 0.8975 761.875 1.3125 ;
      RECT  762.29 0.8975 764.735 1.3125 ;
      RECT  765.15 0.8975 767.595 1.3125 ;
      RECT  768.01 0.8975 770.455 1.3125 ;
      RECT  770.87 0.8975 773.315 1.3125 ;
      RECT  773.73 0.8975 776.175 1.3125 ;
      RECT  776.59 0.8975 779.035 1.3125 ;
      RECT  779.45 0.8975 781.895 1.3125 ;
      RECT  782.31 0.8975 784.755 1.3125 ;
      RECT  785.17 0.8975 787.615 1.3125 ;
      RECT  788.03 0.8975 790.475 1.3125 ;
      RECT  790.89 0.8975 793.335 1.3125 ;
      RECT  793.75 0.8975 796.195 1.3125 ;
      RECT  796.61 0.8975 799.055 1.3125 ;
      RECT  799.47 0.8975 801.915 1.3125 ;
      RECT  802.33 0.8975 804.775 1.3125 ;
      RECT  805.19 0.8975 807.635 1.3125 ;
      RECT  808.05 0.8975 810.495 1.3125 ;
      RECT  810.91 0.8975 813.355 1.3125 ;
      RECT  813.77 0.8975 816.215 1.3125 ;
      RECT  816.63 0.8975 819.075 1.3125 ;
      RECT  819.49 0.8975 821.935 1.3125 ;
      RECT  822.35 0.8975 824.795 1.3125 ;
      RECT  825.21 0.8975 827.655 1.3125 ;
      RECT  828.07 0.8975 830.515 1.3125 ;
      RECT  830.93 0.8975 833.375 1.3125 ;
      RECT  833.79 0.8975 836.235 1.3125 ;
      RECT  836.65 0.8975 839.095 1.3125 ;
      RECT  839.51 0.8975 841.955 1.3125 ;
      RECT  842.37 0.8975 844.815 1.3125 ;
      RECT  845.23 0.8975 847.675 1.3125 ;
      RECT  848.09 0.8975 850.535 1.3125 ;
      RECT  850.95 0.8975 853.395 1.3125 ;
      RECT  853.81 0.8975 856.255 1.3125 ;
      RECT  856.67 0.8975 859.115 1.3125 ;
      RECT  859.53 0.8975 861.975 1.3125 ;
      RECT  862.39 0.8975 864.835 1.3125 ;
      RECT  865.25 0.8975 867.695 1.3125 ;
      RECT  868.11 0.8975 870.555 1.3125 ;
      RECT  870.97 0.8975 873.415 1.3125 ;
      RECT  873.83 0.8975 876.275 1.3125 ;
      RECT  876.69 0.8975 879.135 1.3125 ;
      RECT  879.55 0.8975 881.995 1.3125 ;
      RECT  882.41 0.8975 884.855 1.3125 ;
      RECT  885.27 0.8975 887.715 1.3125 ;
      RECT  888.13 0.8975 890.575 1.3125 ;
      RECT  890.99 0.8975 893.22 1.3125 ;
      RECT  0.14 97.03 64.035 97.445 ;
      RECT  0.14 97.445 64.035 124.97 ;
      RECT  64.035 1.3125 64.45 97.03 ;
      RECT  64.45 97.03 161.275 97.445 ;
      RECT  64.45 97.445 161.275 124.97 ;
      RECT  64.035 97.445 64.45 99.76 ;
      RECT  64.035 100.175 64.45 101.97 ;
      RECT  64.035 102.385 64.45 104.7 ;
      RECT  64.035 105.115 64.45 124.97 ;
      RECT  0.14 1.3125 0.145 60.5 ;
      RECT  0.14 60.5 0.145 60.915 ;
      RECT  0.14 60.915 0.145 97.03 ;
      RECT  0.145 1.3125 0.56 60.5 ;
      RECT  0.56 1.3125 64.035 60.5 ;
      RECT  0.145 60.915 0.56 63.23 ;
      RECT  0.145 63.645 0.56 97.03 ;
      RECT  0.56 60.5 6.3875 60.585 ;
      RECT  0.56 60.585 6.3875 60.915 ;
      RECT  6.3875 60.5 6.8025 60.585 ;
      RECT  6.8025 60.5 64.035 60.585 ;
      RECT  6.8025 60.585 64.035 60.915 ;
      RECT  0.56 60.915 6.3875 61.0 ;
      RECT  0.56 61.0 6.3875 97.03 ;
      RECT  6.3875 61.0 6.8025 97.03 ;
      RECT  6.8025 60.915 64.035 61.0 ;
      RECT  6.8025 61.0 64.035 97.03 ;
      RECT  0.14 0.8975 69.755 1.3125 ;
      RECT  70.17 0.8975 72.615 1.3125 ;
      RECT  73.03 0.8975 75.475 1.3125 ;
      RECT  75.89 0.8975 78.335 1.3125 ;
      RECT  78.75 0.8975 81.195 1.3125 ;
      RECT  81.61 0.8975 84.055 1.3125 ;
      RECT  84.47 0.8975 86.915 1.3125 ;
      RECT  87.33 0.8975 89.775 1.3125 ;
      RECT  90.19 0.8975 92.635 1.3125 ;
      RECT  93.05 0.8975 95.495 1.3125 ;
      RECT  95.91 0.8975 98.355 1.3125 ;
      RECT  98.77 0.8975 101.215 1.3125 ;
      RECT  101.63 0.8975 104.075 1.3125 ;
      RECT  104.49 0.8975 106.935 1.3125 ;
      RECT  107.35 0.8975 109.795 1.3125 ;
      RECT  110.21 0.8975 112.655 1.3125 ;
      RECT  113.07 0.8975 115.515 1.3125 ;
      RECT  115.93 0.8975 118.375 1.3125 ;
      RECT  118.79 0.8975 121.235 1.3125 ;
      RECT  121.65 0.8975 124.095 1.3125 ;
      RECT  124.51 0.8975 126.955 1.3125 ;
      RECT  127.37 0.8975 129.815 1.3125 ;
      RECT  130.23 0.8975 132.675 1.3125 ;
      RECT  133.09 0.8975 135.535 1.3125 ;
      RECT  135.95 0.8975 138.395 1.3125 ;
      RECT  138.81 0.8975 141.255 1.3125 ;
      RECT  141.67 0.8975 144.115 1.3125 ;
      RECT  144.53 0.8975 146.975 1.3125 ;
      RECT  147.39 0.8975 149.835 1.3125 ;
      RECT  150.25 0.8975 152.695 1.3125 ;
      RECT  153.11 0.8975 155.555 1.3125 ;
      RECT  155.97 0.8975 158.415 1.3125 ;
      RECT  158.83 0.8975 161.275 1.3125 ;
      RECT  64.45 1.3125 92.405 71.6425 ;
      RECT  64.45 71.6425 92.405 72.0575 ;
      RECT  64.45 72.0575 92.405 97.03 ;
      RECT  92.405 1.3125 92.82 71.6425 ;
      RECT  92.405 72.0575 92.82 97.03 ;
      RECT  92.82 1.3125 161.275 71.6425 ;
      RECT  92.82 72.0575 161.275 97.03 ;
      RECT  92.82 71.6425 93.11 72.0575 ;
      RECT  93.525 71.6425 93.815 72.0575 ;
      RECT  94.23 71.6425 94.52 72.0575 ;
      RECT  94.935 71.6425 95.225 72.0575 ;
      RECT  95.64 71.6425 95.93 72.0575 ;
      RECT  96.345 71.6425 96.635 72.0575 ;
      RECT  97.05 71.6425 97.34 72.0575 ;
      RECT  97.755 71.6425 98.045 72.0575 ;
      RECT  98.46 71.6425 98.75 72.0575 ;
      RECT  99.165 71.6425 99.455 72.0575 ;
      RECT  99.87 71.6425 100.16 72.0575 ;
      RECT  100.575 71.6425 100.865 72.0575 ;
      RECT  101.28 71.6425 101.57 72.0575 ;
      RECT  101.985 71.6425 102.275 72.0575 ;
      RECT  102.69 71.6425 102.98 72.0575 ;
      RECT  103.395 71.6425 103.685 72.0575 ;
      RECT  104.1 71.6425 104.39 72.0575 ;
      RECT  104.805 71.6425 105.095 72.0575 ;
      RECT  105.51 71.6425 105.8 72.0575 ;
      RECT  106.215 71.6425 106.505 72.0575 ;
      RECT  106.92 71.6425 107.21 72.0575 ;
      RECT  107.625 71.6425 107.915 72.0575 ;
      RECT  108.33 71.6425 108.62 72.0575 ;
      RECT  109.035 71.6425 109.325 72.0575 ;
      RECT  109.74 71.6425 110.03 72.0575 ;
      RECT  110.445 71.6425 110.735 72.0575 ;
      RECT  111.15 71.6425 111.44 72.0575 ;
      RECT  111.855 71.6425 112.145 72.0575 ;
      RECT  112.56 71.6425 112.85 72.0575 ;
      RECT  113.265 71.6425 113.555 72.0575 ;
      RECT  113.97 71.6425 114.26 72.0575 ;
      RECT  114.675 71.6425 114.965 72.0575 ;
      RECT  115.38 71.6425 115.67 72.0575 ;
      RECT  116.085 71.6425 116.375 72.0575 ;
      RECT  116.79 71.6425 117.08 72.0575 ;
      RECT  117.495 71.6425 117.785 72.0575 ;
      RECT  118.2 71.6425 118.49 72.0575 ;
      RECT  118.905 71.6425 119.195 72.0575 ;
      RECT  119.61 71.6425 119.9 72.0575 ;
      RECT  120.315 71.6425 120.605 72.0575 ;
      RECT  121.02 71.6425 121.31 72.0575 ;
      RECT  121.725 71.6425 122.015 72.0575 ;
      RECT  122.43 71.6425 122.72 72.0575 ;
      RECT  123.135 71.6425 123.425 72.0575 ;
      RECT  123.84 71.6425 124.13 72.0575 ;
      RECT  124.545 71.6425 124.835 72.0575 ;
      RECT  125.25 71.6425 125.54 72.0575 ;
      RECT  125.955 71.6425 126.245 72.0575 ;
      RECT  126.66 71.6425 126.95 72.0575 ;
      RECT  127.365 71.6425 127.655 72.0575 ;
      RECT  128.07 71.6425 128.36 72.0575 ;
      RECT  128.775 71.6425 129.065 72.0575 ;
      RECT  129.48 71.6425 129.77 72.0575 ;
      RECT  130.185 71.6425 130.475 72.0575 ;
      RECT  130.89 71.6425 131.18 72.0575 ;
      RECT  131.595 71.6425 131.885 72.0575 ;
      RECT  132.3 71.6425 132.59 72.0575 ;
      RECT  133.005 71.6425 133.295 72.0575 ;
      RECT  133.71 71.6425 134.0 72.0575 ;
      RECT  134.415 71.6425 134.705 72.0575 ;
      RECT  135.12 71.6425 135.41 72.0575 ;
      RECT  135.825 71.6425 136.115 72.0575 ;
      RECT  136.53 71.6425 136.82 72.0575 ;
      RECT  137.235 71.6425 137.525 72.0575 ;
      RECT  137.94 71.6425 138.23 72.0575 ;
      RECT  138.645 71.6425 138.935 72.0575 ;
      RECT  139.35 71.6425 139.64 72.0575 ;
      RECT  140.055 71.6425 140.345 72.0575 ;
      RECT  140.76 71.6425 141.05 72.0575 ;
      RECT  141.465 71.6425 141.755 72.0575 ;
      RECT  142.17 71.6425 142.46 72.0575 ;
      RECT  142.875 71.6425 143.165 72.0575 ;
      RECT  143.58 71.6425 143.87 72.0575 ;
      RECT  144.285 71.6425 144.575 72.0575 ;
      RECT  144.99 71.6425 145.28 72.0575 ;
      RECT  145.695 71.6425 145.985 72.0575 ;
      RECT  146.4 71.6425 146.69 72.0575 ;
      RECT  147.105 71.6425 147.395 72.0575 ;
      RECT  147.81 71.6425 148.1 72.0575 ;
      RECT  148.515 71.6425 148.805 72.0575 ;
      RECT  149.22 71.6425 149.51 72.0575 ;
      RECT  149.925 71.6425 150.215 72.0575 ;
      RECT  150.63 71.6425 150.92 72.0575 ;
      RECT  151.335 71.6425 151.625 72.0575 ;
      RECT  152.04 71.6425 152.33 72.0575 ;
      RECT  152.745 71.6425 153.035 72.0575 ;
      RECT  153.45 71.6425 153.74 72.0575 ;
      RECT  154.155 71.6425 154.445 72.0575 ;
      RECT  154.86 71.6425 155.15 72.0575 ;
      RECT  155.565 71.6425 155.855 72.0575 ;
      RECT  156.27 71.6425 156.56 72.0575 ;
      RECT  156.975 71.6425 157.265 72.0575 ;
      RECT  157.68 71.6425 157.97 72.0575 ;
      RECT  158.385 71.6425 158.675 72.0575 ;
      RECT  159.09 71.6425 159.38 72.0575 ;
      RECT  159.795 71.6425 160.085 72.0575 ;
      RECT  160.5 71.6425 160.79 72.0575 ;
      RECT  161.205 71.6425 161.275 72.0575 ;
      RECT  161.275 1.3125 161.495 71.6425 ;
      RECT  161.275 71.6425 161.495 72.0575 ;
      RECT  161.275 72.0575 161.495 124.97 ;
      RECT  161.495 1.3125 161.69 71.6425 ;
      RECT  161.495 72.0575 161.69 124.97 ;
      RECT  161.69 1.3125 161.91 71.6425 ;
      RECT  161.69 72.0575 161.91 124.97 ;
      RECT  161.91 1.3125 893.22 71.6425 ;
      RECT  161.91 72.0575 893.22 124.97 ;
      RECT  161.91 71.6425 162.2 72.0575 ;
      RECT  162.615 71.6425 162.905 72.0575 ;
      RECT  163.32 71.6425 163.61 72.0575 ;
      RECT  164.025 71.6425 164.315 72.0575 ;
      RECT  164.73 71.6425 165.02 72.0575 ;
      RECT  165.435 71.6425 165.725 72.0575 ;
      RECT  166.14 71.6425 166.43 72.0575 ;
      RECT  166.845 71.6425 167.135 72.0575 ;
      RECT  167.55 71.6425 167.84 72.0575 ;
      RECT  168.255 71.6425 168.545 72.0575 ;
      RECT  168.96 71.6425 169.25 72.0575 ;
      RECT  169.665 71.6425 169.955 72.0575 ;
      RECT  170.37 71.6425 170.66 72.0575 ;
      RECT  171.075 71.6425 171.365 72.0575 ;
      RECT  171.78 71.6425 172.07 72.0575 ;
      RECT  172.485 71.6425 172.775 72.0575 ;
      RECT  173.19 71.6425 173.48 72.0575 ;
      RECT  173.895 71.6425 174.185 72.0575 ;
      RECT  174.6 71.6425 174.89 72.0575 ;
      RECT  175.305 71.6425 175.595 72.0575 ;
      RECT  176.01 71.6425 176.3 72.0575 ;
      RECT  176.715 71.6425 177.005 72.0575 ;
      RECT  177.42 71.6425 177.71 72.0575 ;
      RECT  178.125 71.6425 178.415 72.0575 ;
      RECT  178.83 71.6425 179.12 72.0575 ;
      RECT  179.535 71.6425 179.825 72.0575 ;
      RECT  180.24 71.6425 180.53 72.0575 ;
      RECT  180.945 71.6425 181.235 72.0575 ;
      RECT  181.65 71.6425 181.94 72.0575 ;
      RECT  182.355 71.6425 182.645 72.0575 ;
      RECT  183.06 71.6425 183.35 72.0575 ;
      RECT  183.765 71.6425 184.055 72.0575 ;
      RECT  184.47 71.6425 184.76 72.0575 ;
      RECT  185.175 71.6425 185.465 72.0575 ;
      RECT  185.88 71.6425 186.17 72.0575 ;
      RECT  186.585 71.6425 186.875 72.0575 ;
      RECT  187.29 71.6425 187.58 72.0575 ;
      RECT  187.995 71.6425 188.285 72.0575 ;
      RECT  188.7 71.6425 188.99 72.0575 ;
      RECT  189.405 71.6425 189.695 72.0575 ;
      RECT  190.11 71.6425 190.4 72.0575 ;
      RECT  190.815 71.6425 191.105 72.0575 ;
      RECT  191.52 71.6425 191.81 72.0575 ;
      RECT  192.225 71.6425 192.515 72.0575 ;
      RECT  192.93 71.6425 193.22 72.0575 ;
      RECT  193.635 71.6425 193.925 72.0575 ;
      RECT  194.34 71.6425 194.63 72.0575 ;
      RECT  195.045 71.6425 195.335 72.0575 ;
      RECT  195.75 71.6425 196.04 72.0575 ;
      RECT  196.455 71.6425 196.745 72.0575 ;
      RECT  197.16 71.6425 197.45 72.0575 ;
      RECT  197.865 71.6425 198.155 72.0575 ;
      RECT  198.57 71.6425 198.86 72.0575 ;
      RECT  199.275 71.6425 199.565 72.0575 ;
      RECT  199.98 71.6425 200.27 72.0575 ;
      RECT  200.685 71.6425 200.975 72.0575 ;
      RECT  201.39 71.6425 201.68 72.0575 ;
      RECT  202.095 71.6425 202.385 72.0575 ;
      RECT  202.8 71.6425 203.09 72.0575 ;
      RECT  203.505 71.6425 203.795 72.0575 ;
      RECT  204.21 71.6425 204.5 72.0575 ;
      RECT  204.915 71.6425 205.205 72.0575 ;
      RECT  205.62 71.6425 205.91 72.0575 ;
      RECT  206.325 71.6425 206.615 72.0575 ;
      RECT  207.03 71.6425 207.32 72.0575 ;
      RECT  207.735 71.6425 208.025 72.0575 ;
      RECT  208.44 71.6425 208.73 72.0575 ;
      RECT  209.145 71.6425 209.435 72.0575 ;
      RECT  209.85 71.6425 210.14 72.0575 ;
      RECT  210.555 71.6425 210.845 72.0575 ;
      RECT  211.26 71.6425 211.55 72.0575 ;
      RECT  211.965 71.6425 212.255 72.0575 ;
      RECT  212.67 71.6425 212.96 72.0575 ;
      RECT  213.375 71.6425 213.665 72.0575 ;
      RECT  214.08 71.6425 214.37 72.0575 ;
      RECT  214.785 71.6425 215.075 72.0575 ;
      RECT  215.49 71.6425 215.78 72.0575 ;
      RECT  216.195 71.6425 216.485 72.0575 ;
      RECT  216.9 71.6425 217.19 72.0575 ;
      RECT  217.605 71.6425 217.895 72.0575 ;
      RECT  218.31 71.6425 218.6 72.0575 ;
      RECT  219.015 71.6425 219.305 72.0575 ;
      RECT  219.72 71.6425 220.01 72.0575 ;
      RECT  220.425 71.6425 220.715 72.0575 ;
      RECT  221.13 71.6425 221.42 72.0575 ;
      RECT  221.835 71.6425 222.125 72.0575 ;
      RECT  222.54 71.6425 222.83 72.0575 ;
      RECT  223.245 71.6425 223.535 72.0575 ;
      RECT  223.95 71.6425 224.24 72.0575 ;
      RECT  224.655 71.6425 224.945 72.0575 ;
      RECT  225.36 71.6425 225.65 72.0575 ;
      RECT  226.065 71.6425 226.355 72.0575 ;
      RECT  226.77 71.6425 227.06 72.0575 ;
      RECT  227.475 71.6425 227.765 72.0575 ;
      RECT  228.18 71.6425 228.47 72.0575 ;
      RECT  228.885 71.6425 229.175 72.0575 ;
      RECT  229.59 71.6425 229.88 72.0575 ;
      RECT  230.295 71.6425 230.585 72.0575 ;
      RECT  231.0 71.6425 231.29 72.0575 ;
      RECT  231.705 71.6425 231.995 72.0575 ;
      RECT  232.41 71.6425 232.7 72.0575 ;
      RECT  233.115 71.6425 233.405 72.0575 ;
      RECT  233.82 71.6425 234.11 72.0575 ;
      RECT  234.525 71.6425 234.815 72.0575 ;
      RECT  235.23 71.6425 235.52 72.0575 ;
      RECT  235.935 71.6425 236.225 72.0575 ;
      RECT  236.64 71.6425 236.93 72.0575 ;
      RECT  237.345 71.6425 237.635 72.0575 ;
      RECT  238.05 71.6425 238.34 72.0575 ;
      RECT  238.755 71.6425 239.045 72.0575 ;
      RECT  239.46 71.6425 239.75 72.0575 ;
      RECT  240.165 71.6425 240.455 72.0575 ;
      RECT  240.87 71.6425 241.16 72.0575 ;
      RECT  241.575 71.6425 241.865 72.0575 ;
      RECT  242.28 71.6425 242.57 72.0575 ;
      RECT  242.985 71.6425 243.275 72.0575 ;
      RECT  243.69 71.6425 243.98 72.0575 ;
      RECT  244.395 71.6425 244.685 72.0575 ;
      RECT  245.1 71.6425 245.39 72.0575 ;
      RECT  245.805 71.6425 246.095 72.0575 ;
      RECT  246.51 71.6425 246.8 72.0575 ;
      RECT  247.215 71.6425 247.505 72.0575 ;
      RECT  247.92 71.6425 248.21 72.0575 ;
      RECT  248.625 71.6425 248.915 72.0575 ;
      RECT  249.33 71.6425 249.62 72.0575 ;
      RECT  250.035 71.6425 250.325 72.0575 ;
      RECT  250.74 71.6425 251.03 72.0575 ;
      RECT  251.445 71.6425 251.735 72.0575 ;
      RECT  252.15 71.6425 252.44 72.0575 ;
      RECT  252.855 71.6425 253.145 72.0575 ;
      RECT  253.56 71.6425 253.85 72.0575 ;
      RECT  254.265 71.6425 254.555 72.0575 ;
      RECT  254.97 71.6425 255.26 72.0575 ;
      RECT  255.675 71.6425 255.965 72.0575 ;
      RECT  256.38 71.6425 256.67 72.0575 ;
      RECT  257.085 71.6425 257.375 72.0575 ;
      RECT  257.79 71.6425 258.08 72.0575 ;
      RECT  258.495 71.6425 258.785 72.0575 ;
      RECT  259.2 71.6425 259.49 72.0575 ;
      RECT  259.905 71.6425 260.195 72.0575 ;
      RECT  260.61 71.6425 260.9 72.0575 ;
      RECT  261.315 71.6425 261.605 72.0575 ;
      RECT  262.02 71.6425 262.31 72.0575 ;
      RECT  262.725 71.6425 263.015 72.0575 ;
      RECT  263.43 71.6425 263.72 72.0575 ;
      RECT  264.135 71.6425 264.425 72.0575 ;
      RECT  264.84 71.6425 265.13 72.0575 ;
      RECT  265.545 71.6425 265.835 72.0575 ;
      RECT  266.25 71.6425 266.54 72.0575 ;
      RECT  266.955 71.6425 267.245 72.0575 ;
      RECT  267.66 71.6425 267.95 72.0575 ;
      RECT  268.365 71.6425 268.655 72.0575 ;
      RECT  269.07 71.6425 269.36 72.0575 ;
      RECT  269.775 71.6425 270.065 72.0575 ;
      RECT  270.48 71.6425 270.77 72.0575 ;
      RECT  271.185 71.6425 271.475 72.0575 ;
      RECT  271.89 71.6425 272.18 72.0575 ;
      RECT  272.595 71.6425 893.22 72.0575 ;
   LAYER  metal4 ;
      RECT  0.14 0.14 893.22 124.97 ;
   END
END    mp3_data_array
END    LIBRARY
