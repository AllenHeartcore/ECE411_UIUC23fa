VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO mp3_tag_array_2
   CLASS BLOCK ;
   SIZE 87.995 BY 48.055 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  22.43 1.0375 22.565 1.1725 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  25.29 1.0375 25.425 1.1725 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  28.15 1.0375 28.285 1.1725 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  31.01 1.0375 31.145 1.1725 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  33.87 1.0375 34.005 1.1725 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.73 1.0375 36.865 1.1725 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  39.59 1.0375 39.725 1.1725 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  42.45 1.0375 42.585 1.1725 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.31 1.0375 45.445 1.1725 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  48.17 1.0375 48.305 1.1725 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  51.03 1.0375 51.165 1.1725 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  53.89 1.0375 54.025 1.1725 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.75 1.0375 56.885 1.1725 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.61 1.0375 59.745 1.1725 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  62.47 1.0375 62.605 1.1725 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  65.33 1.0375 65.465 1.1725 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  68.19 1.0375 68.325 1.1725 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.05 1.0375 71.185 1.1725 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.91 1.0375 74.045 1.1725 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.77 1.0375 76.905 1.1725 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  79.63 1.0375 79.765 1.1725 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.49 1.0375 82.625 1.1725 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.35 1.0375 85.485 1.1725 ;
      END
   END din0[22]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  19.57 1.0375 19.705 1.1725 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.85 39.2125 13.985 39.3475 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.85 41.9425 13.985 42.0775 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.85 44.1525 13.985 44.2875 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.85 46.8825 13.985 47.0175 ;
      END
   END addr0[4]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 2.6825 0.42 2.8175 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 5.4125 0.42 5.5475 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.5275 2.7675 6.6625 2.9025 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  31.77 10.87 31.905 11.005 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  33.18 10.87 33.315 11.005 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  34.59 10.87 34.725 11.005 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.0 10.87 36.135 11.005 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.41 10.87 37.545 11.005 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  38.82 10.87 38.955 11.005 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.23 10.87 40.365 11.005 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  41.64 10.87 41.775 11.005 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.05 10.87 43.185 11.005 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  44.46 10.87 44.595 11.005 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.87 10.87 46.005 11.005 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.28 10.87 47.415 11.005 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  48.69 10.87 48.825 11.005 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  50.1 10.87 50.235 11.005 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  51.51 10.87 51.645 11.005 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  52.92 10.87 53.055 11.005 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  54.33 10.87 54.465 11.005 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  55.74 10.87 55.875 11.005 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.15 10.87 57.285 11.005 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  58.56 10.87 58.695 11.005 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.97 10.87 60.105 11.005 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.38 10.87 61.515 11.005 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  62.79 10.87 62.925 11.005 ;
      END
   END dout0[22]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 87.855 47.915 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 87.855 47.915 ;
   LAYER  metal3 ;
      RECT  0.14 0.14 22.29 0.8975 ;
      RECT  22.29 0.14 22.705 0.8975 ;
      RECT  22.29 1.3125 22.705 47.915 ;
      RECT  22.705 0.14 87.855 0.8975 ;
      RECT  22.705 0.8975 25.15 1.3125 ;
      RECT  25.565 0.8975 28.01 1.3125 ;
      RECT  28.425 0.8975 30.87 1.3125 ;
      RECT  31.285 0.8975 33.73 1.3125 ;
      RECT  34.145 0.8975 36.59 1.3125 ;
      RECT  37.005 0.8975 39.45 1.3125 ;
      RECT  39.865 0.8975 42.31 1.3125 ;
      RECT  42.725 0.8975 45.17 1.3125 ;
      RECT  45.585 0.8975 48.03 1.3125 ;
      RECT  48.445 0.8975 50.89 1.3125 ;
      RECT  51.305 0.8975 53.75 1.3125 ;
      RECT  54.165 0.8975 56.61 1.3125 ;
      RECT  57.025 0.8975 59.47 1.3125 ;
      RECT  59.885 0.8975 62.33 1.3125 ;
      RECT  62.745 0.8975 65.19 1.3125 ;
      RECT  65.605 0.8975 68.05 1.3125 ;
      RECT  68.465 0.8975 70.91 1.3125 ;
      RECT  71.325 0.8975 73.77 1.3125 ;
      RECT  74.185 0.8975 76.63 1.3125 ;
      RECT  77.045 0.8975 79.49 1.3125 ;
      RECT  79.905 0.8975 82.35 1.3125 ;
      RECT  82.765 0.8975 85.21 1.3125 ;
      RECT  85.625 0.8975 87.855 1.3125 ;
      RECT  0.14 0.8975 19.43 1.3125 ;
      RECT  19.845 0.8975 22.29 1.3125 ;
      RECT  0.14 39.0725 13.71 39.4875 ;
      RECT  0.14 39.4875 13.71 47.915 ;
      RECT  13.71 1.3125 14.125 39.0725 ;
      RECT  14.125 1.3125 22.29 39.0725 ;
      RECT  14.125 39.0725 22.29 39.4875 ;
      RECT  14.125 39.4875 22.29 47.915 ;
      RECT  13.71 39.4875 14.125 41.8025 ;
      RECT  13.71 42.2175 14.125 44.0125 ;
      RECT  13.71 44.4275 14.125 46.7425 ;
      RECT  13.71 47.1575 14.125 47.915 ;
      RECT  0.14 1.3125 0.145 2.5425 ;
      RECT  0.14 2.5425 0.145 2.9575 ;
      RECT  0.14 2.9575 0.145 39.0725 ;
      RECT  0.145 1.3125 0.56 2.5425 ;
      RECT  0.56 1.3125 13.71 2.5425 ;
      RECT  0.145 2.9575 0.56 5.2725 ;
      RECT  0.145 5.6875 0.56 39.0725 ;
      RECT  0.56 2.5425 6.3875 2.6275 ;
      RECT  0.56 2.6275 6.3875 2.9575 ;
      RECT  6.3875 2.5425 6.8025 2.6275 ;
      RECT  6.8025 2.5425 13.71 2.6275 ;
      RECT  6.8025 2.6275 13.71 2.9575 ;
      RECT  0.56 2.9575 6.3875 3.0425 ;
      RECT  0.56 3.0425 6.3875 39.0725 ;
      RECT  6.3875 3.0425 6.8025 39.0725 ;
      RECT  6.8025 2.9575 13.71 3.0425 ;
      RECT  6.8025 3.0425 13.71 39.0725 ;
      RECT  22.705 1.3125 31.63 10.73 ;
      RECT  22.705 10.73 31.63 11.145 ;
      RECT  22.705 11.145 31.63 47.915 ;
      RECT  31.63 1.3125 32.045 10.73 ;
      RECT  31.63 11.145 32.045 47.915 ;
      RECT  32.045 1.3125 87.855 10.73 ;
      RECT  32.045 11.145 87.855 47.915 ;
      RECT  32.045 10.73 33.04 11.145 ;
      RECT  33.455 10.73 34.45 11.145 ;
      RECT  34.865 10.73 35.86 11.145 ;
      RECT  36.275 10.73 37.27 11.145 ;
      RECT  37.685 10.73 38.68 11.145 ;
      RECT  39.095 10.73 40.09 11.145 ;
      RECT  40.505 10.73 41.5 11.145 ;
      RECT  41.915 10.73 42.91 11.145 ;
      RECT  43.325 10.73 44.32 11.145 ;
      RECT  44.735 10.73 45.73 11.145 ;
      RECT  46.145 10.73 47.14 11.145 ;
      RECT  47.555 10.73 48.55 11.145 ;
      RECT  48.965 10.73 49.96 11.145 ;
      RECT  50.375 10.73 51.37 11.145 ;
      RECT  51.785 10.73 52.78 11.145 ;
      RECT  53.195 10.73 54.19 11.145 ;
      RECT  54.605 10.73 55.6 11.145 ;
      RECT  56.015 10.73 57.01 11.145 ;
      RECT  57.425 10.73 58.42 11.145 ;
      RECT  58.835 10.73 59.83 11.145 ;
      RECT  60.245 10.73 61.24 11.145 ;
      RECT  61.655 10.73 62.65 11.145 ;
      RECT  63.065 10.73 87.855 11.145 ;
   LAYER  metal4 ;
      RECT  0.14 0.14 87.855 47.915 ;
   END
END    mp3_tag_array_2
END    LIBRARY
