VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO mp3_data_array_2
   CLASS BLOCK ;
   SIZE 454.845 BY 96.645 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.98 1.0375 89.115 1.1725 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.84 1.0375 91.975 1.1725 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.7 1.0375 94.835 1.1725 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.56 1.0375 97.695 1.1725 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.42 1.0375 100.555 1.1725 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.28 1.0375 103.415 1.1725 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.14 1.0375 106.275 1.1725 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.0 1.0375 109.135 1.1725 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.86 1.0375 111.995 1.1725 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.72 1.0375 114.855 1.1725 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  117.58 1.0375 117.715 1.1725 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.44 1.0375 120.575 1.1725 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.3 1.0375 123.435 1.1725 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.16 1.0375 126.295 1.1725 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.02 1.0375 129.155 1.1725 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.88 1.0375 132.015 1.1725 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.74 1.0375 134.875 1.1725 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.6 1.0375 137.735 1.1725 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.46 1.0375 140.595 1.1725 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.32 1.0375 143.455 1.1725 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.18 1.0375 146.315 1.1725 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.04 1.0375 149.175 1.1725 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  151.9 1.0375 152.035 1.1725 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  154.76 1.0375 154.895 1.1725 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  157.62 1.0375 157.755 1.1725 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  160.48 1.0375 160.615 1.1725 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  163.34 1.0375 163.475 1.1725 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  166.2 1.0375 166.335 1.1725 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  169.06 1.0375 169.195 1.1725 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  171.92 1.0375 172.055 1.1725 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  174.78 1.0375 174.915 1.1725 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  177.64 1.0375 177.775 1.1725 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  180.5 1.0375 180.635 1.1725 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  183.36 1.0375 183.495 1.1725 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  186.22 1.0375 186.355 1.1725 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  189.08 1.0375 189.215 1.1725 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  191.94 1.0375 192.075 1.1725 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  194.8 1.0375 194.935 1.1725 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  197.66 1.0375 197.795 1.1725 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  200.52 1.0375 200.655 1.1725 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  203.38 1.0375 203.515 1.1725 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  206.24 1.0375 206.375 1.1725 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  209.1 1.0375 209.235 1.1725 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  211.96 1.0375 212.095 1.1725 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  214.82 1.0375 214.955 1.1725 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  217.68 1.0375 217.815 1.1725 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  220.54 1.0375 220.675 1.1725 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  223.4 1.0375 223.535 1.1725 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  226.26 1.0375 226.395 1.1725 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  229.12 1.0375 229.255 1.1725 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  231.98 1.0375 232.115 1.1725 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  234.84 1.0375 234.975 1.1725 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  237.7 1.0375 237.835 1.1725 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  240.56 1.0375 240.695 1.1725 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  243.42 1.0375 243.555 1.1725 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  246.28 1.0375 246.415 1.1725 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  249.14 1.0375 249.275 1.1725 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  252.0 1.0375 252.135 1.1725 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  254.86 1.0375 254.995 1.1725 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  257.72 1.0375 257.855 1.1725 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  260.58 1.0375 260.715 1.1725 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  263.44 1.0375 263.575 1.1725 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  266.3 1.0375 266.435 1.1725 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  269.16 1.0375 269.295 1.1725 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  272.02 1.0375 272.155 1.1725 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  274.88 1.0375 275.015 1.1725 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  277.74 1.0375 277.875 1.1725 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  280.6 1.0375 280.735 1.1725 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  283.46 1.0375 283.595 1.1725 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  286.32 1.0375 286.455 1.1725 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  289.18 1.0375 289.315 1.1725 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  292.04 1.0375 292.175 1.1725 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  294.9 1.0375 295.035 1.1725 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  297.76 1.0375 297.895 1.1725 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  300.62 1.0375 300.755 1.1725 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  303.48 1.0375 303.615 1.1725 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  306.34 1.0375 306.475 1.1725 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  309.2 1.0375 309.335 1.1725 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  312.06 1.0375 312.195 1.1725 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  314.92 1.0375 315.055 1.1725 ;
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  317.78 1.0375 317.915 1.1725 ;
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  320.64 1.0375 320.775 1.1725 ;
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  323.5 1.0375 323.635 1.1725 ;
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  326.36 1.0375 326.495 1.1725 ;
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  329.22 1.0375 329.355 1.1725 ;
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  332.08 1.0375 332.215 1.1725 ;
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  334.94 1.0375 335.075 1.1725 ;
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  337.8 1.0375 337.935 1.1725 ;
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  340.66 1.0375 340.795 1.1725 ;
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  343.52 1.0375 343.655 1.1725 ;
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  346.38 1.0375 346.515 1.1725 ;
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  349.24 1.0375 349.375 1.1725 ;
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  352.1 1.0375 352.235 1.1725 ;
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  354.96 1.0375 355.095 1.1725 ;
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  357.82 1.0375 357.955 1.1725 ;
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  360.68 1.0375 360.815 1.1725 ;
      END
   END din0[95]
   PIN din0[96]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  363.54 1.0375 363.675 1.1725 ;
      END
   END din0[96]
   PIN din0[97]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  366.4 1.0375 366.535 1.1725 ;
      END
   END din0[97]
   PIN din0[98]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  369.26 1.0375 369.395 1.1725 ;
      END
   END din0[98]
   PIN din0[99]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  372.12 1.0375 372.255 1.1725 ;
      END
   END din0[99]
   PIN din0[100]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  374.98 1.0375 375.115 1.1725 ;
      END
   END din0[100]
   PIN din0[101]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  377.84 1.0375 377.975 1.1725 ;
      END
   END din0[101]
   PIN din0[102]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  380.7 1.0375 380.835 1.1725 ;
      END
   END din0[102]
   PIN din0[103]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  383.56 1.0375 383.695 1.1725 ;
      END
   END din0[103]
   PIN din0[104]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  386.42 1.0375 386.555 1.1725 ;
      END
   END din0[104]
   PIN din0[105]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  389.28 1.0375 389.415 1.1725 ;
      END
   END din0[105]
   PIN din0[106]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  392.14 1.0375 392.275 1.1725 ;
      END
   END din0[106]
   PIN din0[107]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  395.0 1.0375 395.135 1.1725 ;
      END
   END din0[107]
   PIN din0[108]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  397.86 1.0375 397.995 1.1725 ;
      END
   END din0[108]
   PIN din0[109]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  400.72 1.0375 400.855 1.1725 ;
      END
   END din0[109]
   PIN din0[110]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  403.58 1.0375 403.715 1.1725 ;
      END
   END din0[110]
   PIN din0[111]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  406.44 1.0375 406.575 1.1725 ;
      END
   END din0[111]
   PIN din0[112]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  409.3 1.0375 409.435 1.1725 ;
      END
   END din0[112]
   PIN din0[113]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  412.16 1.0375 412.295 1.1725 ;
      END
   END din0[113]
   PIN din0[114]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  415.02 1.0375 415.155 1.1725 ;
      END
   END din0[114]
   PIN din0[115]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  417.88 1.0375 418.015 1.1725 ;
      END
   END din0[115]
   PIN din0[116]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  420.74 1.0375 420.875 1.1725 ;
      END
   END din0[116]
   PIN din0[117]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  423.6 1.0375 423.735 1.1725 ;
      END
   END din0[117]
   PIN din0[118]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  426.46 1.0375 426.595 1.1725 ;
      END
   END din0[118]
   PIN din0[119]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  429.32 1.0375 429.455 1.1725 ;
      END
   END din0[119]
   PIN din0[120]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  432.18 1.0375 432.315 1.1725 ;
      END
   END din0[120]
   PIN din0[121]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  435.04 1.0375 435.175 1.1725 ;
      END
   END din0[121]
   PIN din0[122]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  437.9 1.0375 438.035 1.1725 ;
      END
   END din0[122]
   PIN din0[123]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  440.76 1.0375 440.895 1.1725 ;
      END
   END din0[123]
   PIN din0[124]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  443.62 1.0375 443.755 1.1725 ;
      END
   END din0[124]
   PIN din0[125]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  446.48 1.0375 446.615 1.1725 ;
      END
   END din0[125]
   PIN din0[126]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  449.34 1.0375 449.475 1.1725 ;
      END
   END din0[126]
   PIN din0[127]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  452.2 1.0375 452.335 1.1725 ;
      END
   END din0[127]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.5 71.55 37.635 71.685 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.5 74.28 37.635 74.415 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.5 76.49 37.635 76.625 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.5 79.22 37.635 79.355 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.5 81.43 37.635 81.565 ;
      END
   END addr0[4]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 29.56 0.42 29.695 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 32.29 0.42 32.425 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.5275 29.645 6.6625 29.78 ;
      END
   END clk0
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.22 1.0375 43.355 1.1725 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  46.08 1.0375 46.215 1.1725 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  48.94 1.0375 49.075 1.1725 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  51.8 1.0375 51.935 1.1725 ;
      END
   END wmask0[3]
   PIN wmask0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  54.66 1.0375 54.795 1.1725 ;
      END
   END wmask0[4]
   PIN wmask0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  57.52 1.0375 57.655 1.1725 ;
      END
   END wmask0[5]
   PIN wmask0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.38 1.0375 60.515 1.1725 ;
      END
   END wmask0[6]
   PIN wmask0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.24 1.0375 63.375 1.1725 ;
      END
   END wmask0[7]
   PIN wmask0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.1 1.0375 66.235 1.1725 ;
      END
   END wmask0[8]
   PIN wmask0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  68.96 1.0375 69.095 1.1725 ;
      END
   END wmask0[9]
   PIN wmask0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.82 1.0375 71.955 1.1725 ;
      END
   END wmask0[10]
   PIN wmask0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  74.68 1.0375 74.815 1.1725 ;
      END
   END wmask0[11]
   PIN wmask0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  77.54 1.0375 77.675 1.1725 ;
      END
   END wmask0[12]
   PIN wmask0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.4 1.0375 80.535 1.1725 ;
      END
   END wmask0[13]
   PIN wmask0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.26 1.0375 83.395 1.1725 ;
      END
   END wmask0[14]
   PIN wmask0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.12 1.0375 86.255 1.1725 ;
      END
   END wmask0[15]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.01 40.7025 61.145 40.8375 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.715 40.7025 61.85 40.8375 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  62.42 40.7025 62.555 40.8375 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.125 40.7025 63.26 40.8375 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  63.83 40.7025 63.965 40.8375 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.535 40.7025 64.67 40.8375 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  65.24 40.7025 65.375 40.8375 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  65.945 40.7025 66.08 40.8375 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  66.65 40.7025 66.785 40.8375 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.355 40.7025 67.49 40.8375 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  68.06 40.7025 68.195 40.8375 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  68.765 40.7025 68.9 40.8375 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  69.47 40.7025 69.605 40.8375 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.175 40.7025 70.31 40.8375 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.88 40.7025 71.015 40.8375 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  71.585 40.7025 71.72 40.8375 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.29 40.7025 72.425 40.8375 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  72.995 40.7025 73.13 40.8375 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.7 40.7025 73.835 40.8375 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  74.405 40.7025 74.54 40.8375 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.11 40.7025 75.245 40.8375 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  75.815 40.7025 75.95 40.8375 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.52 40.7025 76.655 40.8375 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  77.225 40.7025 77.36 40.8375 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  77.93 40.7025 78.065 40.8375 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  78.635 40.7025 78.77 40.8375 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  79.34 40.7025 79.475 40.8375 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.045 40.7025 80.18 40.8375 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  80.75 40.7025 80.885 40.8375 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.455 40.7025 81.59 40.8375 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.16 40.7025 82.295 40.8375 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  82.865 40.7025 83.0 40.8375 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  83.57 40.7025 83.705 40.8375 ;
      END
   END dout0[32]
   PIN dout0[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  84.275 40.7025 84.41 40.8375 ;
      END
   END dout0[33]
   PIN dout0[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  84.98 40.7025 85.115 40.8375 ;
      END
   END dout0[34]
   PIN dout0[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  85.685 40.7025 85.82 40.8375 ;
      END
   END dout0[35]
   PIN dout0[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  86.39 40.7025 86.525 40.8375 ;
      END
   END dout0[36]
   PIN dout0[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  87.095 40.7025 87.23 40.8375 ;
      END
   END dout0[37]
   PIN dout0[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  87.8 40.7025 87.935 40.8375 ;
      END
   END dout0[38]
   PIN dout0[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  88.505 40.7025 88.64 40.8375 ;
      END
   END dout0[39]
   PIN dout0[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.21 40.7025 89.345 40.8375 ;
      END
   END dout0[40]
   PIN dout0[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  89.915 40.7025 90.05 40.8375 ;
      END
   END dout0[41]
   PIN dout0[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  90.62 40.7025 90.755 40.8375 ;
      END
   END dout0[42]
   PIN dout0[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  91.325 40.7025 91.46 40.8375 ;
      END
   END dout0[43]
   PIN dout0[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.03 40.7025 92.165 40.8375 ;
      END
   END dout0[44]
   PIN dout0[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  92.735 40.7025 92.87 40.8375 ;
      END
   END dout0[45]
   PIN dout0[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  93.44 40.7025 93.575 40.8375 ;
      END
   END dout0[46]
   PIN dout0[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.145 40.7025 94.28 40.8375 ;
      END
   END dout0[47]
   PIN dout0[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  94.85 40.7025 94.985 40.8375 ;
      END
   END dout0[48]
   PIN dout0[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  95.555 40.7025 95.69 40.8375 ;
      END
   END dout0[49]
   PIN dout0[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.26 40.7025 96.395 40.8375 ;
      END
   END dout0[50]
   PIN dout0[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  96.965 40.7025 97.1 40.8375 ;
      END
   END dout0[51]
   PIN dout0[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  97.67 40.7025 97.805 40.8375 ;
      END
   END dout0[52]
   PIN dout0[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  98.375 40.7025 98.51 40.8375 ;
      END
   END dout0[53]
   PIN dout0[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.08 40.7025 99.215 40.8375 ;
      END
   END dout0[54]
   PIN dout0[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  99.785 40.7025 99.92 40.8375 ;
      END
   END dout0[55]
   PIN dout0[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  100.49 40.7025 100.625 40.8375 ;
      END
   END dout0[56]
   PIN dout0[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.195 40.7025 101.33 40.8375 ;
      END
   END dout0[57]
   PIN dout0[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  101.9 40.7025 102.035 40.8375 ;
      END
   END dout0[58]
   PIN dout0[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  102.605 40.7025 102.74 40.8375 ;
      END
   END dout0[59]
   PIN dout0[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  103.31 40.7025 103.445 40.8375 ;
      END
   END dout0[60]
   PIN dout0[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.015 40.7025 104.15 40.8375 ;
      END
   END dout0[61]
   PIN dout0[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  104.72 40.7025 104.855 40.8375 ;
      END
   END dout0[62]
   PIN dout0[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  105.425 40.7025 105.56 40.8375 ;
      END
   END dout0[63]
   PIN dout0[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.13 40.7025 106.265 40.8375 ;
      END
   END dout0[64]
   PIN dout0[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  106.835 40.7025 106.97 40.8375 ;
      END
   END dout0[65]
   PIN dout0[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  107.54 40.7025 107.675 40.8375 ;
      END
   END dout0[66]
   PIN dout0[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.245 40.7025 108.38 40.8375 ;
      END
   END dout0[67]
   PIN dout0[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  108.95 40.7025 109.085 40.8375 ;
      END
   END dout0[68]
   PIN dout0[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  109.655 40.7025 109.79 40.8375 ;
      END
   END dout0[69]
   PIN dout0[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  110.36 40.7025 110.495 40.8375 ;
      END
   END dout0[70]
   PIN dout0[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.065 40.7025 111.2 40.8375 ;
      END
   END dout0[71]
   PIN dout0[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  111.77 40.7025 111.905 40.8375 ;
      END
   END dout0[72]
   PIN dout0[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  112.475 40.7025 112.61 40.8375 ;
      END
   END dout0[73]
   PIN dout0[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.18 40.7025 113.315 40.8375 ;
      END
   END dout0[74]
   PIN dout0[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  113.885 40.7025 114.02 40.8375 ;
      END
   END dout0[75]
   PIN dout0[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  114.59 40.7025 114.725 40.8375 ;
      END
   END dout0[76]
   PIN dout0[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  115.295 40.7025 115.43 40.8375 ;
      END
   END dout0[77]
   PIN dout0[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  116.0 40.7025 116.135 40.8375 ;
      END
   END dout0[78]
   PIN dout0[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  116.705 40.7025 116.84 40.8375 ;
      END
   END dout0[79]
   PIN dout0[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  117.41 40.7025 117.545 40.8375 ;
      END
   END dout0[80]
   PIN dout0[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.115 40.7025 118.25 40.8375 ;
      END
   END dout0[81]
   PIN dout0[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  118.82 40.7025 118.955 40.8375 ;
      END
   END dout0[82]
   PIN dout0[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  119.525 40.7025 119.66 40.8375 ;
      END
   END dout0[83]
   PIN dout0[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.23 40.7025 120.365 40.8375 ;
      END
   END dout0[84]
   PIN dout0[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  120.935 40.7025 121.07 40.8375 ;
      END
   END dout0[85]
   PIN dout0[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  121.64 40.7025 121.775 40.8375 ;
      END
   END dout0[86]
   PIN dout0[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  122.345 40.7025 122.48 40.8375 ;
      END
   END dout0[87]
   PIN dout0[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.05 40.7025 123.185 40.8375 ;
      END
   END dout0[88]
   PIN dout0[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  123.755 40.7025 123.89 40.8375 ;
      END
   END dout0[89]
   PIN dout0[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  124.46 40.7025 124.595 40.8375 ;
      END
   END dout0[90]
   PIN dout0[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  125.165 40.7025 125.3 40.8375 ;
      END
   END dout0[91]
   PIN dout0[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  125.87 40.7025 126.005 40.8375 ;
      END
   END dout0[92]
   PIN dout0[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  126.575 40.7025 126.71 40.8375 ;
      END
   END dout0[93]
   PIN dout0[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  127.28 40.7025 127.415 40.8375 ;
      END
   END dout0[94]
   PIN dout0[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  127.985 40.7025 128.12 40.8375 ;
      END
   END dout0[95]
   PIN dout0[96]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  128.69 40.7025 128.825 40.8375 ;
      END
   END dout0[96]
   PIN dout0[97]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  129.395 40.7025 129.53 40.8375 ;
      END
   END dout0[97]
   PIN dout0[98]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  130.1 40.7025 130.235 40.8375 ;
      END
   END dout0[98]
   PIN dout0[99]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  130.805 40.7025 130.94 40.8375 ;
      END
   END dout0[99]
   PIN dout0[100]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  131.51 40.7025 131.645 40.8375 ;
      END
   END dout0[100]
   PIN dout0[101]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.215 40.7025 132.35 40.8375 ;
      END
   END dout0[101]
   PIN dout0[102]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  132.92 40.7025 133.055 40.8375 ;
      END
   END dout0[102]
   PIN dout0[103]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  133.625 40.7025 133.76 40.8375 ;
      END
   END dout0[103]
   PIN dout0[104]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  134.33 40.7025 134.465 40.8375 ;
      END
   END dout0[104]
   PIN dout0[105]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.035 40.7025 135.17 40.8375 ;
      END
   END dout0[105]
   PIN dout0[106]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  135.74 40.7025 135.875 40.8375 ;
      END
   END dout0[106]
   PIN dout0[107]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  136.445 40.7025 136.58 40.8375 ;
      END
   END dout0[107]
   PIN dout0[108]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.15 40.7025 137.285 40.8375 ;
      END
   END dout0[108]
   PIN dout0[109]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.855 40.7025 137.99 40.8375 ;
      END
   END dout0[109]
   PIN dout0[110]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  138.56 40.7025 138.695 40.8375 ;
      END
   END dout0[110]
   PIN dout0[111]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  139.265 40.7025 139.4 40.8375 ;
      END
   END dout0[111]
   PIN dout0[112]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  139.97 40.7025 140.105 40.8375 ;
      END
   END dout0[112]
   PIN dout0[113]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  140.675 40.7025 140.81 40.8375 ;
      END
   END dout0[113]
   PIN dout0[114]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  141.38 40.7025 141.515 40.8375 ;
      END
   END dout0[114]
   PIN dout0[115]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  142.085 40.7025 142.22 40.8375 ;
      END
   END dout0[115]
   PIN dout0[116]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  142.79 40.7025 142.925 40.8375 ;
      END
   END dout0[116]
   PIN dout0[117]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  143.495 40.7025 143.63 40.8375 ;
      END
   END dout0[117]
   PIN dout0[118]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  144.2 40.7025 144.335 40.8375 ;
      END
   END dout0[118]
   PIN dout0[119]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  144.905 40.7025 145.04 40.8375 ;
      END
   END dout0[119]
   PIN dout0[120]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  145.61 40.7025 145.745 40.8375 ;
      END
   END dout0[120]
   PIN dout0[121]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  146.315 40.7025 146.45 40.8375 ;
      END
   END dout0[121]
   PIN dout0[122]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  147.02 40.7025 147.155 40.8375 ;
      END
   END dout0[122]
   PIN dout0[123]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  147.725 40.7025 147.86 40.8375 ;
      END
   END dout0[123]
   PIN dout0[124]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  148.43 40.7025 148.565 40.8375 ;
      END
   END dout0[124]
   PIN dout0[125]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.135 40.7025 149.27 40.8375 ;
      END
   END dout0[125]
   PIN dout0[126]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  149.84 40.7025 149.975 40.8375 ;
      END
   END dout0[126]
   PIN dout0[127]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  150.545 40.7025 150.68 40.8375 ;
      END
   END dout0[127]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 454.705 96.505 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 454.705 96.505 ;
   LAYER  metal3 ;
      RECT  0.14 0.14 88.84 0.8975 ;
      RECT  88.84 0.14 89.255 0.8975 ;
      RECT  89.255 0.14 454.705 0.8975 ;
      RECT  89.255 0.8975 91.7 1.3125 ;
      RECT  92.115 0.8975 94.56 1.3125 ;
      RECT  94.975 0.8975 97.42 1.3125 ;
      RECT  97.835 0.8975 100.28 1.3125 ;
      RECT  100.695 0.8975 103.14 1.3125 ;
      RECT  103.555 0.8975 106.0 1.3125 ;
      RECT  106.415 0.8975 108.86 1.3125 ;
      RECT  109.275 0.8975 111.72 1.3125 ;
      RECT  112.135 0.8975 114.58 1.3125 ;
      RECT  114.995 0.8975 117.44 1.3125 ;
      RECT  117.855 0.8975 120.3 1.3125 ;
      RECT  120.715 0.8975 123.16 1.3125 ;
      RECT  123.575 0.8975 126.02 1.3125 ;
      RECT  126.435 0.8975 128.88 1.3125 ;
      RECT  129.295 0.8975 131.74 1.3125 ;
      RECT  132.155 0.8975 134.6 1.3125 ;
      RECT  135.015 0.8975 137.46 1.3125 ;
      RECT  137.875 0.8975 140.32 1.3125 ;
      RECT  140.735 0.8975 143.18 1.3125 ;
      RECT  143.595 0.8975 146.04 1.3125 ;
      RECT  146.455 0.8975 148.9 1.3125 ;
      RECT  149.315 0.8975 151.76 1.3125 ;
      RECT  152.175 0.8975 154.62 1.3125 ;
      RECT  155.035 0.8975 157.48 1.3125 ;
      RECT  157.895 0.8975 160.34 1.3125 ;
      RECT  160.755 0.8975 163.2 1.3125 ;
      RECT  163.615 0.8975 166.06 1.3125 ;
      RECT  166.475 0.8975 168.92 1.3125 ;
      RECT  169.335 0.8975 171.78 1.3125 ;
      RECT  172.195 0.8975 174.64 1.3125 ;
      RECT  175.055 0.8975 177.5 1.3125 ;
      RECT  177.915 0.8975 180.36 1.3125 ;
      RECT  180.775 0.8975 183.22 1.3125 ;
      RECT  183.635 0.8975 186.08 1.3125 ;
      RECT  186.495 0.8975 188.94 1.3125 ;
      RECT  189.355 0.8975 191.8 1.3125 ;
      RECT  192.215 0.8975 194.66 1.3125 ;
      RECT  195.075 0.8975 197.52 1.3125 ;
      RECT  197.935 0.8975 200.38 1.3125 ;
      RECT  200.795 0.8975 203.24 1.3125 ;
      RECT  203.655 0.8975 206.1 1.3125 ;
      RECT  206.515 0.8975 208.96 1.3125 ;
      RECT  209.375 0.8975 211.82 1.3125 ;
      RECT  212.235 0.8975 214.68 1.3125 ;
      RECT  215.095 0.8975 217.54 1.3125 ;
      RECT  217.955 0.8975 220.4 1.3125 ;
      RECT  220.815 0.8975 223.26 1.3125 ;
      RECT  223.675 0.8975 226.12 1.3125 ;
      RECT  226.535 0.8975 228.98 1.3125 ;
      RECT  229.395 0.8975 231.84 1.3125 ;
      RECT  232.255 0.8975 234.7 1.3125 ;
      RECT  235.115 0.8975 237.56 1.3125 ;
      RECT  237.975 0.8975 240.42 1.3125 ;
      RECT  240.835 0.8975 243.28 1.3125 ;
      RECT  243.695 0.8975 246.14 1.3125 ;
      RECT  246.555 0.8975 249.0 1.3125 ;
      RECT  249.415 0.8975 251.86 1.3125 ;
      RECT  252.275 0.8975 254.72 1.3125 ;
      RECT  255.135 0.8975 257.58 1.3125 ;
      RECT  257.995 0.8975 260.44 1.3125 ;
      RECT  260.855 0.8975 263.3 1.3125 ;
      RECT  263.715 0.8975 266.16 1.3125 ;
      RECT  266.575 0.8975 269.02 1.3125 ;
      RECT  269.435 0.8975 271.88 1.3125 ;
      RECT  272.295 0.8975 274.74 1.3125 ;
      RECT  275.155 0.8975 277.6 1.3125 ;
      RECT  278.015 0.8975 280.46 1.3125 ;
      RECT  280.875 0.8975 283.32 1.3125 ;
      RECT  283.735 0.8975 286.18 1.3125 ;
      RECT  286.595 0.8975 289.04 1.3125 ;
      RECT  289.455 0.8975 291.9 1.3125 ;
      RECT  292.315 0.8975 294.76 1.3125 ;
      RECT  295.175 0.8975 297.62 1.3125 ;
      RECT  298.035 0.8975 300.48 1.3125 ;
      RECT  300.895 0.8975 303.34 1.3125 ;
      RECT  303.755 0.8975 306.2 1.3125 ;
      RECT  306.615 0.8975 309.06 1.3125 ;
      RECT  309.475 0.8975 311.92 1.3125 ;
      RECT  312.335 0.8975 314.78 1.3125 ;
      RECT  315.195 0.8975 317.64 1.3125 ;
      RECT  318.055 0.8975 320.5 1.3125 ;
      RECT  320.915 0.8975 323.36 1.3125 ;
      RECT  323.775 0.8975 326.22 1.3125 ;
      RECT  326.635 0.8975 329.08 1.3125 ;
      RECT  329.495 0.8975 331.94 1.3125 ;
      RECT  332.355 0.8975 334.8 1.3125 ;
      RECT  335.215 0.8975 337.66 1.3125 ;
      RECT  338.075 0.8975 340.52 1.3125 ;
      RECT  340.935 0.8975 343.38 1.3125 ;
      RECT  343.795 0.8975 346.24 1.3125 ;
      RECT  346.655 0.8975 349.1 1.3125 ;
      RECT  349.515 0.8975 351.96 1.3125 ;
      RECT  352.375 0.8975 354.82 1.3125 ;
      RECT  355.235 0.8975 357.68 1.3125 ;
      RECT  358.095 0.8975 360.54 1.3125 ;
      RECT  360.955 0.8975 363.4 1.3125 ;
      RECT  363.815 0.8975 366.26 1.3125 ;
      RECT  366.675 0.8975 369.12 1.3125 ;
      RECT  369.535 0.8975 371.98 1.3125 ;
      RECT  372.395 0.8975 374.84 1.3125 ;
      RECT  375.255 0.8975 377.7 1.3125 ;
      RECT  378.115 0.8975 380.56 1.3125 ;
      RECT  380.975 0.8975 383.42 1.3125 ;
      RECT  383.835 0.8975 386.28 1.3125 ;
      RECT  386.695 0.8975 389.14 1.3125 ;
      RECT  389.555 0.8975 392.0 1.3125 ;
      RECT  392.415 0.8975 394.86 1.3125 ;
      RECT  395.275 0.8975 397.72 1.3125 ;
      RECT  398.135 0.8975 400.58 1.3125 ;
      RECT  400.995 0.8975 403.44 1.3125 ;
      RECT  403.855 0.8975 406.3 1.3125 ;
      RECT  406.715 0.8975 409.16 1.3125 ;
      RECT  409.575 0.8975 412.02 1.3125 ;
      RECT  412.435 0.8975 414.88 1.3125 ;
      RECT  415.295 0.8975 417.74 1.3125 ;
      RECT  418.155 0.8975 420.6 1.3125 ;
      RECT  421.015 0.8975 423.46 1.3125 ;
      RECT  423.875 0.8975 426.32 1.3125 ;
      RECT  426.735 0.8975 429.18 1.3125 ;
      RECT  429.595 0.8975 432.04 1.3125 ;
      RECT  432.455 0.8975 434.9 1.3125 ;
      RECT  435.315 0.8975 437.76 1.3125 ;
      RECT  438.175 0.8975 440.62 1.3125 ;
      RECT  441.035 0.8975 443.48 1.3125 ;
      RECT  443.895 0.8975 446.34 1.3125 ;
      RECT  446.755 0.8975 449.2 1.3125 ;
      RECT  449.615 0.8975 452.06 1.3125 ;
      RECT  452.475 0.8975 454.705 1.3125 ;
      RECT  0.14 71.41 37.36 71.825 ;
      RECT  0.14 71.825 37.36 96.505 ;
      RECT  37.36 1.3125 37.775 71.41 ;
      RECT  37.775 71.41 88.84 71.825 ;
      RECT  37.775 71.825 88.84 96.505 ;
      RECT  37.36 71.825 37.775 74.14 ;
      RECT  37.36 74.555 37.775 76.35 ;
      RECT  37.36 76.765 37.775 79.08 ;
      RECT  37.36 79.495 37.775 81.29 ;
      RECT  37.36 81.705 37.775 96.505 ;
      RECT  0.14 1.3125 0.145 29.42 ;
      RECT  0.14 29.42 0.145 29.835 ;
      RECT  0.14 29.835 0.145 71.41 ;
      RECT  0.145 1.3125 0.56 29.42 ;
      RECT  0.56 1.3125 37.36 29.42 ;
      RECT  0.145 29.835 0.56 32.15 ;
      RECT  0.145 32.565 0.56 71.41 ;
      RECT  0.56 29.42 6.3875 29.505 ;
      RECT  0.56 29.505 6.3875 29.835 ;
      RECT  6.3875 29.42 6.8025 29.505 ;
      RECT  6.8025 29.42 37.36 29.505 ;
      RECT  6.8025 29.505 37.36 29.835 ;
      RECT  0.56 29.835 6.3875 29.92 ;
      RECT  0.56 29.92 6.3875 71.41 ;
      RECT  6.3875 29.92 6.8025 71.41 ;
      RECT  6.8025 29.835 37.36 29.92 ;
      RECT  6.8025 29.92 37.36 71.41 ;
      RECT  0.14 0.8975 43.08 1.3125 ;
      RECT  43.495 0.8975 45.94 1.3125 ;
      RECT  46.355 0.8975 48.8 1.3125 ;
      RECT  49.215 0.8975 51.66 1.3125 ;
      RECT  52.075 0.8975 54.52 1.3125 ;
      RECT  54.935 0.8975 57.38 1.3125 ;
      RECT  57.795 0.8975 60.24 1.3125 ;
      RECT  60.655 0.8975 63.1 1.3125 ;
      RECT  63.515 0.8975 65.96 1.3125 ;
      RECT  66.375 0.8975 68.82 1.3125 ;
      RECT  69.235 0.8975 71.68 1.3125 ;
      RECT  72.095 0.8975 74.54 1.3125 ;
      RECT  74.955 0.8975 77.4 1.3125 ;
      RECT  77.815 0.8975 80.26 1.3125 ;
      RECT  80.675 0.8975 83.12 1.3125 ;
      RECT  83.535 0.8975 85.98 1.3125 ;
      RECT  86.395 0.8975 88.84 1.3125 ;
      RECT  37.775 1.3125 60.87 40.5625 ;
      RECT  37.775 40.5625 60.87 40.9775 ;
      RECT  37.775 40.9775 60.87 71.41 ;
      RECT  60.87 1.3125 61.285 40.5625 ;
      RECT  60.87 40.9775 61.285 71.41 ;
      RECT  61.285 1.3125 88.84 40.5625 ;
      RECT  61.285 40.9775 88.84 71.41 ;
      RECT  61.285 40.5625 61.575 40.9775 ;
      RECT  61.99 40.5625 62.28 40.9775 ;
      RECT  62.695 40.5625 62.985 40.9775 ;
      RECT  63.4 40.5625 63.69 40.9775 ;
      RECT  64.105 40.5625 64.395 40.9775 ;
      RECT  64.81 40.5625 65.1 40.9775 ;
      RECT  65.515 40.5625 65.805 40.9775 ;
      RECT  66.22 40.5625 66.51 40.9775 ;
      RECT  66.925 40.5625 67.215 40.9775 ;
      RECT  67.63 40.5625 67.92 40.9775 ;
      RECT  68.335 40.5625 68.625 40.9775 ;
      RECT  69.04 40.5625 69.33 40.9775 ;
      RECT  69.745 40.5625 70.035 40.9775 ;
      RECT  70.45 40.5625 70.74 40.9775 ;
      RECT  71.155 40.5625 71.445 40.9775 ;
      RECT  71.86 40.5625 72.15 40.9775 ;
      RECT  72.565 40.5625 72.855 40.9775 ;
      RECT  73.27 40.5625 73.56 40.9775 ;
      RECT  73.975 40.5625 74.265 40.9775 ;
      RECT  74.68 40.5625 74.97 40.9775 ;
      RECT  75.385 40.5625 75.675 40.9775 ;
      RECT  76.09 40.5625 76.38 40.9775 ;
      RECT  76.795 40.5625 77.085 40.9775 ;
      RECT  77.5 40.5625 77.79 40.9775 ;
      RECT  78.205 40.5625 78.495 40.9775 ;
      RECT  78.91 40.5625 79.2 40.9775 ;
      RECT  79.615 40.5625 79.905 40.9775 ;
      RECT  80.32 40.5625 80.61 40.9775 ;
      RECT  81.025 40.5625 81.315 40.9775 ;
      RECT  81.73 40.5625 82.02 40.9775 ;
      RECT  82.435 40.5625 82.725 40.9775 ;
      RECT  83.14 40.5625 83.43 40.9775 ;
      RECT  83.845 40.5625 84.135 40.9775 ;
      RECT  84.55 40.5625 84.84 40.9775 ;
      RECT  85.255 40.5625 85.545 40.9775 ;
      RECT  85.96 40.5625 86.25 40.9775 ;
      RECT  86.665 40.5625 86.955 40.9775 ;
      RECT  87.37 40.5625 87.66 40.9775 ;
      RECT  88.075 40.5625 88.365 40.9775 ;
      RECT  88.78 40.5625 88.84 40.9775 ;
      RECT  88.84 1.3125 89.07 40.5625 ;
      RECT  88.84 40.5625 89.07 40.9775 ;
      RECT  88.84 40.9775 89.07 96.505 ;
      RECT  89.07 1.3125 89.255 40.5625 ;
      RECT  89.07 40.9775 89.255 96.505 ;
      RECT  89.255 1.3125 89.485 40.5625 ;
      RECT  89.255 40.9775 89.485 96.505 ;
      RECT  89.485 1.3125 454.705 40.5625 ;
      RECT  89.485 40.9775 454.705 96.505 ;
      RECT  89.485 40.5625 89.775 40.9775 ;
      RECT  90.19 40.5625 90.48 40.9775 ;
      RECT  90.895 40.5625 91.185 40.9775 ;
      RECT  91.6 40.5625 91.89 40.9775 ;
      RECT  92.305 40.5625 92.595 40.9775 ;
      RECT  93.01 40.5625 93.3 40.9775 ;
      RECT  93.715 40.5625 94.005 40.9775 ;
      RECT  94.42 40.5625 94.71 40.9775 ;
      RECT  95.125 40.5625 95.415 40.9775 ;
      RECT  95.83 40.5625 96.12 40.9775 ;
      RECT  96.535 40.5625 96.825 40.9775 ;
      RECT  97.24 40.5625 97.53 40.9775 ;
      RECT  97.945 40.5625 98.235 40.9775 ;
      RECT  98.65 40.5625 98.94 40.9775 ;
      RECT  99.355 40.5625 99.645 40.9775 ;
      RECT  100.06 40.5625 100.35 40.9775 ;
      RECT  100.765 40.5625 101.055 40.9775 ;
      RECT  101.47 40.5625 101.76 40.9775 ;
      RECT  102.175 40.5625 102.465 40.9775 ;
      RECT  102.88 40.5625 103.17 40.9775 ;
      RECT  103.585 40.5625 103.875 40.9775 ;
      RECT  104.29 40.5625 104.58 40.9775 ;
      RECT  104.995 40.5625 105.285 40.9775 ;
      RECT  105.7 40.5625 105.99 40.9775 ;
      RECT  106.405 40.5625 106.695 40.9775 ;
      RECT  107.11 40.5625 107.4 40.9775 ;
      RECT  107.815 40.5625 108.105 40.9775 ;
      RECT  108.52 40.5625 108.81 40.9775 ;
      RECT  109.225 40.5625 109.515 40.9775 ;
      RECT  109.93 40.5625 110.22 40.9775 ;
      RECT  110.635 40.5625 110.925 40.9775 ;
      RECT  111.34 40.5625 111.63 40.9775 ;
      RECT  112.045 40.5625 112.335 40.9775 ;
      RECT  112.75 40.5625 113.04 40.9775 ;
      RECT  113.455 40.5625 113.745 40.9775 ;
      RECT  114.16 40.5625 114.45 40.9775 ;
      RECT  114.865 40.5625 115.155 40.9775 ;
      RECT  115.57 40.5625 115.86 40.9775 ;
      RECT  116.275 40.5625 116.565 40.9775 ;
      RECT  116.98 40.5625 117.27 40.9775 ;
      RECT  117.685 40.5625 117.975 40.9775 ;
      RECT  118.39 40.5625 118.68 40.9775 ;
      RECT  119.095 40.5625 119.385 40.9775 ;
      RECT  119.8 40.5625 120.09 40.9775 ;
      RECT  120.505 40.5625 120.795 40.9775 ;
      RECT  121.21 40.5625 121.5 40.9775 ;
      RECT  121.915 40.5625 122.205 40.9775 ;
      RECT  122.62 40.5625 122.91 40.9775 ;
      RECT  123.325 40.5625 123.615 40.9775 ;
      RECT  124.03 40.5625 124.32 40.9775 ;
      RECT  124.735 40.5625 125.025 40.9775 ;
      RECT  125.44 40.5625 125.73 40.9775 ;
      RECT  126.145 40.5625 126.435 40.9775 ;
      RECT  126.85 40.5625 127.14 40.9775 ;
      RECT  127.555 40.5625 127.845 40.9775 ;
      RECT  128.26 40.5625 128.55 40.9775 ;
      RECT  128.965 40.5625 129.255 40.9775 ;
      RECT  129.67 40.5625 129.96 40.9775 ;
      RECT  130.375 40.5625 130.665 40.9775 ;
      RECT  131.08 40.5625 131.37 40.9775 ;
      RECT  131.785 40.5625 132.075 40.9775 ;
      RECT  132.49 40.5625 132.78 40.9775 ;
      RECT  133.195 40.5625 133.485 40.9775 ;
      RECT  133.9 40.5625 134.19 40.9775 ;
      RECT  134.605 40.5625 134.895 40.9775 ;
      RECT  135.31 40.5625 135.6 40.9775 ;
      RECT  136.015 40.5625 136.305 40.9775 ;
      RECT  136.72 40.5625 137.01 40.9775 ;
      RECT  137.425 40.5625 137.715 40.9775 ;
      RECT  138.13 40.5625 138.42 40.9775 ;
      RECT  138.835 40.5625 139.125 40.9775 ;
      RECT  139.54 40.5625 139.83 40.9775 ;
      RECT  140.245 40.5625 140.535 40.9775 ;
      RECT  140.95 40.5625 141.24 40.9775 ;
      RECT  141.655 40.5625 141.945 40.9775 ;
      RECT  142.36 40.5625 142.65 40.9775 ;
      RECT  143.065 40.5625 143.355 40.9775 ;
      RECT  143.77 40.5625 144.06 40.9775 ;
      RECT  144.475 40.5625 144.765 40.9775 ;
      RECT  145.18 40.5625 145.47 40.9775 ;
      RECT  145.885 40.5625 146.175 40.9775 ;
      RECT  146.59 40.5625 146.88 40.9775 ;
      RECT  147.295 40.5625 147.585 40.9775 ;
      RECT  148.0 40.5625 148.29 40.9775 ;
      RECT  148.705 40.5625 148.995 40.9775 ;
      RECT  149.41 40.5625 149.7 40.9775 ;
      RECT  150.115 40.5625 150.405 40.9775 ;
      RECT  150.82 40.5625 454.705 40.9775 ;
   LAYER  metal4 ;
      RECT  0.14 0.14 454.705 96.505 ;
   END
END    mp3_data_array_2
END    LIBRARY
