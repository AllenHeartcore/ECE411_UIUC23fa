module top;
import mult_types::*;

    multiplier_itf itf();
    grader grd (.*);
    testbench tb (.*);
endmodule : top
