VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO mp3_tag_array
   CLASS BLOCK ;
   SIZE 84.585 BY 46.5 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  19.02 1.0375 19.155 1.1725 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  21.88 1.0375 22.015 1.1725 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  24.74 1.0375 24.875 1.1725 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  27.6 1.0375 27.735 1.1725 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  30.46 1.0375 30.595 1.1725 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  33.32 1.0375 33.455 1.1725 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.18 1.0375 36.315 1.1725 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  39.04 1.0375 39.175 1.1725 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  41.9 1.0375 42.035 1.1725 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  44.76 1.0375 44.895 1.1725 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  47.62 1.0375 47.755 1.1725 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  50.48 1.0375 50.615 1.1725 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  53.34 1.0375 53.475 1.1725 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  56.2 1.0375 56.335 1.1725 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  59.06 1.0375 59.195 1.1725 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  61.92 1.0375 62.055 1.1725 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  64.78 1.0375 64.915 1.1725 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.64 1.0375 67.775 1.1725 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  70.5 1.0375 70.635 1.1725 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  73.36 1.0375 73.495 1.1725 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  76.22 1.0375 76.355 1.1725 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  79.08 1.0375 79.215 1.1725 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  81.94 1.0375 82.075 1.1725 ;
      END
   END din0[22]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.3 37.6575 13.435 37.7925 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.3 40.3875 13.435 40.5225 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.3 42.5975 13.435 42.7325 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  13.3 45.3275 13.435 45.4625 ;
      END
   END addr0[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 1.1275 0.42 1.2625 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.285 3.8575 0.42 3.9925 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  6.5275 1.2125 6.6625 1.3475 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  29.845 12.27 29.98 12.405 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  30.55 12.27 30.685 12.405 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  31.255 12.27 31.39 12.405 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  31.96 12.27 32.095 12.405 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.665 12.27 32.8 12.405 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  33.37 12.27 33.505 12.405 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  34.075 12.27 34.21 12.405 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  34.78 12.27 34.915 12.405 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  35.485 12.27 35.62 12.405 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.19 12.27 36.325 12.405 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  36.895 12.27 37.03 12.405 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  37.6 12.27 37.735 12.405 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  38.305 12.27 38.44 12.405 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  39.01 12.27 39.145 12.405 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  39.715 12.27 39.85 12.405 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  40.42 12.27 40.555 12.405 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  41.125 12.27 41.26 12.405 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  41.83 12.27 41.965 12.405 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  42.535 12.27 42.67 12.405 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.24 12.27 43.375 12.405 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  43.945 12.27 44.08 12.405 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  44.65 12.27 44.785 12.405 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  45.355 12.27 45.49 12.405 ;
      END
   END dout0[22]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 84.445 46.36 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 84.445 46.36 ;
   LAYER  metal3 ;
      RECT  0.14 0.14 18.88 0.8975 ;
      RECT  18.88 0.14 19.295 0.8975 ;
      RECT  18.88 1.3125 19.295 46.36 ;
      RECT  19.295 0.14 84.445 0.8975 ;
      RECT  19.295 0.8975 21.74 1.3125 ;
      RECT  22.155 0.8975 24.6 1.3125 ;
      RECT  25.015 0.8975 27.46 1.3125 ;
      RECT  27.875 0.8975 30.32 1.3125 ;
      RECT  30.735 0.8975 33.18 1.3125 ;
      RECT  33.595 0.8975 36.04 1.3125 ;
      RECT  36.455 0.8975 38.9 1.3125 ;
      RECT  39.315 0.8975 41.76 1.3125 ;
      RECT  42.175 0.8975 44.62 1.3125 ;
      RECT  45.035 0.8975 47.48 1.3125 ;
      RECT  47.895 0.8975 50.34 1.3125 ;
      RECT  50.755 0.8975 53.2 1.3125 ;
      RECT  53.615 0.8975 56.06 1.3125 ;
      RECT  56.475 0.8975 58.92 1.3125 ;
      RECT  59.335 0.8975 61.78 1.3125 ;
      RECT  62.195 0.8975 64.64 1.3125 ;
      RECT  65.055 0.8975 67.5 1.3125 ;
      RECT  67.915 0.8975 70.36 1.3125 ;
      RECT  70.775 0.8975 73.22 1.3125 ;
      RECT  73.635 0.8975 76.08 1.3125 ;
      RECT  76.495 0.8975 78.94 1.3125 ;
      RECT  79.355 0.8975 81.8 1.3125 ;
      RECT  82.215 0.8975 84.445 1.3125 ;
      RECT  0.14 37.5175 13.16 37.9325 ;
      RECT  0.14 37.9325 13.16 46.36 ;
      RECT  13.16 1.3125 13.575 37.5175 ;
      RECT  13.575 1.3125 18.88 37.5175 ;
      RECT  13.575 37.5175 18.88 37.9325 ;
      RECT  13.575 37.9325 18.88 46.36 ;
      RECT  13.16 37.9325 13.575 40.2475 ;
      RECT  13.16 40.6625 13.575 42.4575 ;
      RECT  13.16 42.8725 13.575 45.1875 ;
      RECT  13.16 45.6025 13.575 46.36 ;
      RECT  0.14 0.8975 0.145 0.9875 ;
      RECT  0.14 0.9875 0.145 1.3125 ;
      RECT  0.145 0.8975 0.56 0.9875 ;
      RECT  0.56 0.8975 18.88 0.9875 ;
      RECT  0.14 1.3125 0.145 1.4025 ;
      RECT  0.14 1.4025 0.145 37.5175 ;
      RECT  0.145 1.4025 0.56 3.7175 ;
      RECT  0.145 4.1325 0.56 37.5175 ;
      RECT  0.56 0.9875 6.3875 1.0725 ;
      RECT  0.56 1.0725 6.3875 1.3125 ;
      RECT  6.3875 0.9875 6.8025 1.0725 ;
      RECT  6.8025 0.9875 18.88 1.0725 ;
      RECT  6.8025 1.0725 18.88 1.3125 ;
      RECT  0.56 1.3125 6.3875 1.4025 ;
      RECT  6.8025 1.3125 13.16 1.4025 ;
      RECT  0.56 1.4025 6.3875 1.4875 ;
      RECT  0.56 1.4875 6.3875 37.5175 ;
      RECT  6.3875 1.4875 6.8025 37.5175 ;
      RECT  6.8025 1.4025 13.16 1.4875 ;
      RECT  6.8025 1.4875 13.16 37.5175 ;
      RECT  19.295 1.3125 29.705 12.13 ;
      RECT  19.295 12.13 29.705 12.545 ;
      RECT  19.295 12.545 29.705 46.36 ;
      RECT  29.705 1.3125 30.12 12.13 ;
      RECT  29.705 12.545 30.12 46.36 ;
      RECT  30.12 1.3125 84.445 12.13 ;
      RECT  30.12 12.545 84.445 46.36 ;
      RECT  30.12 12.13 30.41 12.545 ;
      RECT  30.825 12.13 31.115 12.545 ;
      RECT  31.53 12.13 31.82 12.545 ;
      RECT  32.235 12.13 32.525 12.545 ;
      RECT  32.94 12.13 33.23 12.545 ;
      RECT  33.645 12.13 33.935 12.545 ;
      RECT  34.35 12.13 34.64 12.545 ;
      RECT  35.055 12.13 35.345 12.545 ;
      RECT  35.76 12.13 36.05 12.545 ;
      RECT  36.465 12.13 36.755 12.545 ;
      RECT  37.17 12.13 37.46 12.545 ;
      RECT  37.875 12.13 38.165 12.545 ;
      RECT  38.58 12.13 38.87 12.545 ;
      RECT  39.285 12.13 39.575 12.545 ;
      RECT  39.99 12.13 40.28 12.545 ;
      RECT  40.695 12.13 40.985 12.545 ;
      RECT  41.4 12.13 41.69 12.545 ;
      RECT  42.105 12.13 42.395 12.545 ;
      RECT  42.81 12.13 43.1 12.545 ;
      RECT  43.515 12.13 43.805 12.545 ;
      RECT  44.22 12.13 44.51 12.545 ;
      RECT  44.925 12.13 45.215 12.545 ;
      RECT  45.63 12.13 84.445 12.545 ;
   LAYER  metal4 ;
      RECT  0.14 0.14 84.445 46.36 ;
   END
END    mp3_tag_array
END    LIBRARY
